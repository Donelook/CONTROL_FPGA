-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 7 2025 00:28:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49287\ : std_logic;
signal \N__49280\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49271\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49260\ : std_logic;
signal \N__49253\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49251\ : std_logic;
signal \N__49244\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49242\ : std_logic;
signal \N__49225\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49213\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49208\ : std_logic;
signal \N__49205\ : std_logic;
signal \N__49202\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49192\ : std_logic;
signal \N__49189\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49183\ : std_logic;
signal \N__49180\ : std_logic;
signal \N__49177\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49165\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49149\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49138\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49124\ : std_logic;
signal \N__49121\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49115\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49111\ : std_logic;
signal \N__49108\ : std_logic;
signal \N__49105\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49103\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49100\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49088\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49069\ : std_logic;
signal \N__49066\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49039\ : std_logic;
signal \N__49036\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49018\ : std_logic;
signal \N__49015\ : std_logic;
signal \N__49014\ : std_logic;
signal \N__49013\ : std_logic;
signal \N__49010\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49002\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48996\ : std_logic;
signal \N__48993\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48973\ : std_logic;
signal \N__48972\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48949\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48925\ : std_logic;
signal \N__48922\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48908\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48871\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48841\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48833\ : std_logic;
signal \N__48832\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48830\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48827\ : std_logic;
signal \N__48826\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48824\ : std_logic;
signal \N__48823\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48820\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48817\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48814\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48811\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48808\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48805\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48802\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48794\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48791\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48788\ : std_logic;
signal \N__48787\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48784\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48778\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48773\ : std_logic;
signal \N__48772\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48770\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48767\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48764\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48761\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48755\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48752\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48747\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48743\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48740\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48735\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48732\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48727\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48721\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48718\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48715\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48712\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48345\ : std_logic;
signal \N__48344\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48312\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48303\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48276\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48233\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48200\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48172\ : std_logic;
signal \N__48171\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48161\ : std_logic;
signal \N__48160\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48155\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48149\ : std_logic;
signal \N__48148\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48146\ : std_logic;
signal \N__48145\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48137\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48134\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48130\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48124\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48122\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48103\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48100\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48097\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48089\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47776\ : std_logic;
signal \N__47773\ : std_logic;
signal \N__47772\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47765\ : std_logic;
signal \N__47762\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47713\ : std_logic;
signal \N__47710\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47704\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47680\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47636\ : std_logic;
signal \N__47633\ : std_logic;
signal \N__47630\ : std_logic;
signal \N__47627\ : std_logic;
signal \N__47622\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47608\ : std_logic;
signal \N__47605\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47600\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47575\ : std_logic;
signal \N__47572\ : std_logic;
signal \N__47569\ : std_logic;
signal \N__47566\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47561\ : std_logic;
signal \N__47558\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47394\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47365\ : std_logic;
signal \N__47364\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47362\ : std_logic;
signal \N__47361\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47351\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47345\ : std_logic;
signal \N__47342\ : std_logic;
signal \N__47339\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47306\ : std_logic;
signal \N__47303\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47293\ : std_logic;
signal \N__47290\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47282\ : std_logic;
signal \N__47279\ : std_logic;
signal \N__47276\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47257\ : std_logic;
signal \N__47254\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47249\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47238\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47228\ : std_logic;
signal \N__47225\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47199\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47192\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47151\ : std_logic;
signal \N__47148\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47139\ : std_logic;
signal \N__47138\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47108\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47102\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47096\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46924\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46899\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46884\ : std_logic;
signal \N__46883\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46877\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46864\ : std_logic;
signal \N__46861\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46856\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46834\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46828\ : std_logic;
signal \N__46825\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46810\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46789\ : std_logic;
signal \N__46788\ : std_logic;
signal \N__46785\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46770\ : std_logic;
signal \N__46765\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46754\ : std_logic;
signal \N__46751\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46709\ : std_logic;
signal \N__46706\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46693\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46669\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46663\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46645\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46642\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46632\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46616\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46610\ : std_logic;
signal \N__46607\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46580\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46486\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46473\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46454\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46427\ : std_logic;
signal \N__46424\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46417\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46415\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46390\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46379\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46361\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46344\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46337\ : std_logic;
signal \N__46334\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46325\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46305\ : std_logic;
signal \N__46302\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46262\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46241\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46235\ : std_logic;
signal \N__46232\ : std_logic;
signal \N__46229\ : std_logic;
signal \N__46226\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46220\ : std_logic;
signal \N__46219\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46184\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46174\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46153\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46135\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46129\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46094\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46048\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46030\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45983\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45973\ : std_logic;
signal \N__45970\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45951\ : std_logic;
signal \N__45948\ : std_logic;
signal \N__45945\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45923\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45893\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45861\ : std_logic;
signal \N__45858\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45852\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45823\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45818\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45802\ : std_logic;
signal \N__45799\ : std_logic;
signal \N__45796\ : std_logic;
signal \N__45793\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45784\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45775\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45771\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45757\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45723\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45713\ : std_logic;
signal \N__45710\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45663\ : std_logic;
signal \N__45660\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45653\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45634\ : std_logic;
signal \N__45631\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45628\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45625\ : std_logic;
signal \N__45622\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45615\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45609\ : std_logic;
signal \N__45604\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45560\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45547\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45512\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45509\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45506\ : std_logic;
signal \N__45505\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45503\ : std_logic;
signal \N__45502\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45500\ : std_logic;
signal \N__45499\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45434\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45386\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45379\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45375\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45366\ : std_logic;
signal \N__45365\ : std_logic;
signal \N__45362\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45320\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45287\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45270\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45264\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45253\ : std_logic;
signal \N__45250\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45226\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45206\ : std_logic;
signal \N__45203\ : std_logic;
signal \N__45200\ : std_logic;
signal \N__45197\ : std_logic;
signal \N__45196\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45166\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45161\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45157\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45154\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45142\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45137\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45131\ : std_logic;
signal \N__45128\ : std_logic;
signal \N__45125\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45119\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45106\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45094\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45006\ : std_logic;
signal \N__45005\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44993\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44975\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44966\ : std_logic;
signal \N__44963\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44913\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44845\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44836\ : std_logic;
signal \N__44833\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44811\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44798\ : std_logic;
signal \N__44795\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44773\ : std_logic;
signal \N__44770\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44760\ : std_logic;
signal \N__44757\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44742\ : std_logic;
signal \N__44737\ : std_logic;
signal \N__44734\ : std_logic;
signal \N__44731\ : std_logic;
signal \N__44728\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44569\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44561\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44559\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44556\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44551\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44526\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44461\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44446\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44390\ : std_logic;
signal \N__44387\ : std_logic;
signal \N__44384\ : std_logic;
signal \N__44377\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44337\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44313\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44302\ : std_logic;
signal \N__44299\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44281\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44215\ : std_logic;
signal \N__44212\ : std_logic;
signal \N__44209\ : std_logic;
signal \N__44206\ : std_logic;
signal \N__44203\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44094\ : std_logic;
signal \N__44091\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44083\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44080\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44059\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44056\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44029\ : std_logic;
signal \N__44026\ : std_logic;
signal \N__44023\ : std_logic;
signal \N__44020\ : std_logic;
signal \N__44017\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44011\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43986\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43970\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43944\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43937\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43921\ : std_logic;
signal \N__43918\ : std_logic;
signal \N__43915\ : std_logic;
signal \N__43912\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43877\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43851\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43840\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43788\ : std_logic;
signal \N__43783\ : std_logic;
signal \N__43780\ : std_logic;
signal \N__43777\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43753\ : std_logic;
signal \N__43750\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43744\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43737\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43714\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43708\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43705\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43694\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43647\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43644\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43531\ : std_logic;
signal \N__43528\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43522\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43516\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43500\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43498\ : std_logic;
signal \N__43497\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43495\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43490\ : std_logic;
signal \N__43483\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43469\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43467\ : std_logic;
signal \N__43466\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43464\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43458\ : std_logic;
signal \N__43457\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43454\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43451\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43434\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43430\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43424\ : std_logic;
signal \N__43421\ : std_logic;
signal \N__43418\ : std_logic;
signal \N__43415\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43394\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43388\ : std_logic;
signal \N__43385\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43364\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43361\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43358\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43350\ : std_logic;
signal \N__43345\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43341\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43338\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43326\ : std_logic;
signal \N__43317\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43301\ : std_logic;
signal \N__43294\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43247\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43223\ : std_logic;
signal \N__43220\ : std_logic;
signal \N__43217\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43187\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43148\ : std_logic;
signal \N__43145\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43057\ : std_logic;
signal \N__43054\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43027\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43019\ : std_logic;
signal \N__43016\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42993\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42978\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42958\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42943\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42929\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42903\ : std_logic;
signal \N__42900\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42810\ : std_logic;
signal \N__42807\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42772\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42764\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42741\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42730\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42700\ : std_logic;
signal \N__42699\ : std_logic;
signal \N__42696\ : std_logic;
signal \N__42693\ : std_logic;
signal \N__42690\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42642\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42630\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42595\ : std_logic;
signal \N__42592\ : std_logic;
signal \N__42591\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42588\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42549\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42535\ : std_logic;
signal \N__42532\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42474\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42438\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42414\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42394\ : std_logic;
signal \N__42391\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42332\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42328\ : std_logic;
signal \N__42325\ : std_logic;
signal \N__42322\ : std_logic;
signal \N__42319\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42317\ : std_logic;
signal \N__42316\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42313\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42308\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42305\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42287\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42270\ : std_logic;
signal \N__42267\ : std_logic;
signal \N__42264\ : std_logic;
signal \N__42261\ : std_logic;
signal \N__42254\ : std_logic;
signal \N__42251\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42237\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42214\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42179\ : std_logic;
signal \N__42178\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42173\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42134\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42080\ : std_logic;
signal \N__42077\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42058\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42056\ : std_logic;
signal \N__42055\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42049\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42003\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41994\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41962\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41956\ : std_logic;
signal \N__41953\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41938\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41908\ : std_logic;
signal \N__41905\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41890\ : std_logic;
signal \N__41887\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41857\ : std_logic;
signal \N__41854\ : std_logic;
signal \N__41851\ : std_logic;
signal \N__41848\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41794\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41779\ : std_logic;
signal \N__41776\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41770\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41764\ : std_logic;
signal \N__41761\ : std_logic;
signal \N__41758\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41750\ : std_logic;
signal \N__41747\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41731\ : std_logic;
signal \N__41728\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41706\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41702\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41686\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41654\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41629\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41590\ : std_logic;
signal \N__41587\ : std_logic;
signal \N__41584\ : std_logic;
signal \N__41581\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41546\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41540\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41520\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41511\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41501\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41447\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41434\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41391\ : std_logic;
signal \N__41388\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41384\ : std_logic;
signal \N__41381\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41358\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41337\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41311\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41287\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41267\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41261\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41207\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41140\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41108\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41102\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41090\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41074\ : std_logic;
signal \N__41071\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41052\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41036\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41015\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40989\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40983\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40959\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40894\ : std_logic;
signal \N__40891\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40867\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40862\ : std_logic;
signal \N__40859\ : std_logic;
signal \N__40856\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40843\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40832\ : std_logic;
signal \N__40829\ : std_logic;
signal \N__40826\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40818\ : std_logic;
signal \N__40815\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40808\ : std_logic;
signal \N__40805\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40793\ : std_logic;
signal \N__40790\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40774\ : std_logic;
signal \N__40771\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40765\ : std_logic;
signal \N__40764\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40749\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40701\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40691\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40673\ : std_logic;
signal \N__40670\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40636\ : std_logic;
signal \N__40633\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40541\ : std_logic;
signal \N__40538\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40532\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40522\ : std_logic;
signal \N__40521\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40499\ : std_logic;
signal \N__40496\ : std_logic;
signal \N__40493\ : std_logic;
signal \N__40490\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40481\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40472\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40463\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40439\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40372\ : std_logic;
signal \N__40369\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40340\ : std_logic;
signal \N__40337\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40313\ : std_logic;
signal \N__40310\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40300\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40295\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40289\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40273\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40259\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40244\ : std_logic;
signal \N__40243\ : std_logic;
signal \N__40240\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40222\ : std_logic;
signal \N__40219\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40211\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40193\ : std_logic;
signal \N__40190\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40184\ : std_logic;
signal \N__40181\ : std_logic;
signal \N__40178\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40118\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40109\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40092\ : std_logic;
signal \N__40089\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40083\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40070\ : std_logic;
signal \N__40065\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40010\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39953\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39947\ : std_logic;
signal \N__39944\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39929\ : std_logic;
signal \N__39926\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39917\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39911\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39898\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39892\ : std_logic;
signal \N__39889\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39883\ : std_logic;
signal \N__39880\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39862\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39821\ : std_logic;
signal \N__39818\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39763\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39755\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39740\ : std_logic;
signal \N__39737\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39691\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39655\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39632\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39553\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39549\ : std_logic;
signal \N__39546\ : std_logic;
signal \N__39545\ : std_logic;
signal \N__39542\ : std_logic;
signal \N__39539\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39466\ : std_logic;
signal \N__39463\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39249\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39235\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39214\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39208\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39181\ : std_logic;
signal \N__39178\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39172\ : std_logic;
signal \N__39169\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39161\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39124\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39091\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39082\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39055\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39046\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38989\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38983\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38974\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38884\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38864\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38810\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38798\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38792\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38722\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38695\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38647\ : std_logic;
signal \N__38644\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38560\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38542\ : std_logic;
signal \N__38539\ : std_logic;
signal \N__38536\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38437\ : std_logic;
signal \N__38434\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38410\ : std_logic;
signal \N__38407\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38338\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38287\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38200\ : std_logic;
signal \N__38197\ : std_logic;
signal \N__38194\ : std_logic;
signal \N__38191\ : std_logic;
signal \N__38188\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37951\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37945\ : std_logic;
signal \N__37942\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37936\ : std_logic;
signal \N__37933\ : std_logic;
signal \N__37930\ : std_logic;
signal \N__37927\ : std_logic;
signal \N__37924\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37918\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37903\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37858\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37849\ : std_logic;
signal \N__37846\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37831\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37816\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37750\ : std_logic;
signal \N__37747\ : std_logic;
signal \N__37744\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37729\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37717\ : std_logic;
signal \N__37714\ : std_logic;
signal \N__37711\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37687\ : std_logic;
signal \N__37684\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37660\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37618\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37561\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37552\ : std_logic;
signal \N__37549\ : std_logic;
signal \N__37546\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37513\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37504\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37489\ : std_logic;
signal \N__37486\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37474\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37450\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37402\ : std_logic;
signal \N__37399\ : std_logic;
signal \N__37394\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37381\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37321\ : std_logic;
signal \N__37318\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37285\ : std_logic;
signal \N__37282\ : std_logic;
signal \N__37277\ : std_logic;
signal \N__37274\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37261\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37246\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37228\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37216\ : std_logic;
signal \N__37213\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37172\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37166\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37142\ : std_logic;
signal \N__37139\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37060\ : std_logic;
signal \N__37057\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37051\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37030\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36989\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36931\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36886\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36853\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36769\ : std_logic;
signal \N__36766\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36757\ : std_logic;
signal \N__36754\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36748\ : std_logic;
signal \N__36745\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36709\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36581\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36541\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36525\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36445\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36442\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36437\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36398\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36316\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36149\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35801\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35737\ : std_logic;
signal \N__35734\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35556\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35349\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35229\ : std_logic;
signal \N__35226\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35108\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34826\ : std_logic;
signal \N__34823\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34580\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34478\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34402\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34324\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34081\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33605\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33593\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33259\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32574\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32146\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32056\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32044\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31846\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31844\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31729\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31714\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31705\ : std_logic;
signal \N__31702\ : std_logic;
signal \N__31699\ : std_logic;
signal \N__31696\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31684\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31657\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31558\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31546\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31531\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31516\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31363\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31328\ : std_logic;
signal \N__31325\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31277\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31210\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30851\ : std_logic;
signal \N__30848\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30806\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30512\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30294\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30263\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30193\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29692\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29554\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29333\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29278\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28317\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27973\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27967\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27274\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25655\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25652\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25532\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25433\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24079\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23931\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21528\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20000\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1_16\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal \current_shift_inst.PI_CTRL.m14_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_19_cascade_\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_7\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_4\ : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_10 : std_logic;
signal \current_shift_inst.PI_CTRL.m7_2\ : std_logic;
signal pwm_duty_input_7 : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_15\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_20\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_8\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_2_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_118\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_178\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \N_22_i_i\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_6\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\ : std_logic;
signal pwm_duty_input_6 : std_logic;
signal i8_mux : std_logic;
signal \N_28_mux\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_0\ : std_logic;
signal \bfn_3_9_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_8\ : std_logic;
signal \bfn_3_10_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_acc_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_3_11_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_acc_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\ : std_logic;
signal \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \clk_10khz_RNIIENAZ0Z2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \bfn_4_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \bfn_4_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal un7_start_stop_0_a3 : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal un5_counter_cry_1 : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal un5_counter_cry_2 : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal un5_counter_cry_3 : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal un5_counter_cry_4 : std_logic;
signal \counterZ0Z_6\ : std_logic;
signal un5_counter_cry_5 : std_logic;
signal \counter_RNO_0Z0Z_7\ : std_logic;
signal un5_counter_cry_6 : std_logic;
signal un5_counter_cry_7 : std_logic;
signal un5_counter_cry_8 : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \counter_RNO_0Z0Z_10\ : std_logic;
signal un5_counter_cry_9 : std_logic;
signal un5_counter_cry_10 : std_logic;
signal un5_counter_cry_11 : std_logic;
signal \counter_RNO_0Z0Z_12\ : std_logic;
signal \counterZ0Z_10\ : std_logic;
signal \counterZ0Z_7\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \un2_counter_5_cascade_\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \counterZ0Z_11\ : std_logic;
signal \counterZ0Z_9\ : std_logic;
signal \counterZ0Z_12\ : std_logic;
signal \counterZ0Z_8\ : std_logic;
signal un2_counter_7 : std_logic;
signal un2_counter_8 : std_logic;
signal un2_counter_9 : std_logic;
signal clk_10khz_i : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_enablelt3_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_0\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_16_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47_21_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_7\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_2\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_3\ : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.N_228_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_0\ : std_logic;
signal \bfn_8_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \bfn_8_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \bfn_8_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.N_199\ : std_logic;
signal \current_shift_inst.phase_validZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3\ : std_logic;
signal measured_delay_hc_21 : std_logic;
signal measured_delay_hc_20 : std_logic;
signal measured_delay_hc_22 : std_logic;
signal \pwm_generator_inst.threshold_ACCZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt15\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \pwm_generator_inst.thresholdZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_75\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_76\ : std_logic;
signal \N_717_g\ : std_logic;
signal \current_shift_inst.meas_stateZ0Z_0\ : std_logic;
signal \current_shift_inst.S3_riseZ0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z0\ : std_logic;
signal \current_shift_inst.S3_syncZ0Z1\ : std_logic;
signal \current_shift_inst.S3_sync_prevZ0\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\ : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal delay_hc_d2 : std_logic;
signal measured_delay_hc_26 : std_logic;
signal measured_delay_hc_30 : std_logic;
signal measured_delay_hc_25 : std_logic;
signal measured_delay_hc_23 : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_29 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto13\ : std_logic;
signal measured_delay_hc_19 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\ : std_logic;
signal \bfn_10_12_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_10_13_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.N_232_cascade_\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_21_cascade_\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \current_shift_inst.z_i_0_31\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_2\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILORI_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_13\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI190J_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_15\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_18\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_21\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\ : std_logic;
signal \bfn_10_24_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_23\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_26\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_27\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_28\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_29\ : std_logic;
signal \current_shift_inst.un38_control_input_0_cry_30\ : std_logic;
signal \bfn_10_25_0_\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_25\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_336_i\ : std_logic;
signal measured_delay_hc_27 : std_logic;
signal measured_delay_hc_28 : std_logic;
signal il_min_comp1_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2_cascade_\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst1.N_231\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \current_shift_inst.S1_riseZ0\ : std_logic;
signal \current_shift_inst.S1_syncZ0Z0\ : std_logic;
signal \phase_controller_inst1.start_timer_tr_0_sqmuxa\ : std_logic;
signal \current_shift_inst.S1_syncZ0Z1\ : std_logic;
signal \current_shift_inst.S1_sync_prevZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_0\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_0\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_1_cry_0\ : std_logic;
signal \current_shift_inst.control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_8\ : std_logic;
signal \bfn_11_21_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_16\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \current_shift_inst.control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.control_inputZ0Z_24\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \current_shift_inst.phase_valid_RNISLORZ0Z2\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24\ : std_logic;
signal \current_shift_inst.control_input_1_cry_24_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_336_i_g\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal s1_phy_c : std_logic;
signal \phase_controller_inst1.stoper_tr.N_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3\ : std_logic;
signal \current_shift_inst.z_i_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_12_24_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \bfn_12_25_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_12_26_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_337_i\ : std_logic;
signal start_stop_c : std_logic;
signal red_c_i : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\ : std_logic;
signal \current_shift_inst.un38_control_input_0_axb_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\ : std_logic;
signal \current_shift_inst.start_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.stop_timer_phaseZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\ : std_logic;
signal \current_shift_inst.timer_phase.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_13_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal s2_phy_c : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto31_0_0\ : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal measured_delay_hc_16 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_18 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_1\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_3\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_fast_31\ : std_logic;
signal \G_407\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\ : std_logic;
signal \G_406\ : std_logic;
signal \current_shift_inst.z_cry_0\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\ : std_logic;
signal \current_shift_inst.z_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\ : std_logic;
signal \current_shift_inst.z_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\ : std_logic;
signal \current_shift_inst.z_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\ : std_logic;
signal \current_shift_inst.z_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\ : std_logic;
signal \current_shift_inst.z_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\ : std_logic;
signal \current_shift_inst.z_cry_6\ : std_logic;
signal \current_shift_inst.z_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\ : std_logic;
signal \current_shift_inst.z_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\ : std_logic;
signal \current_shift_inst.z_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\ : std_logic;
signal \current_shift_inst.z_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\ : std_logic;
signal \current_shift_inst.z_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\ : std_logic;
signal \current_shift_inst.z_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\ : std_logic;
signal \current_shift_inst.z_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\ : std_logic;
signal \current_shift_inst.z_cry_14\ : std_logic;
signal \current_shift_inst.z_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\ : std_logic;
signal \current_shift_inst.z_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\ : std_logic;
signal \current_shift_inst.z_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\ : std_logic;
signal \current_shift_inst.z_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\ : std_logic;
signal \current_shift_inst.z_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\ : std_logic;
signal \current_shift_inst.z_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\ : std_logic;
signal \current_shift_inst.z_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\ : std_logic;
signal \current_shift_inst.z_cry_22\ : std_logic;
signal \current_shift_inst.z_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\ : std_logic;
signal \bfn_14_21_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\ : std_logic;
signal \current_shift_inst.z_cry_24\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\ : std_logic;
signal \current_shift_inst.z_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\ : std_logic;
signal \current_shift_inst.z_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\ : std_logic;
signal \current_shift_inst.z_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\ : std_logic;
signal \current_shift_inst.z_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\ : std_logic;
signal \current_shift_inst.z_cry_29\ : std_logic;
signal \current_shift_inst.z_cry_30\ : std_logic;
signal \current_shift_inst.z_31\ : std_logic;
signal \bfn_14_22_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_7\ : std_logic;
signal \bfn_14_23_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_15\ : std_logic;
signal \bfn_14_24_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_23\ : std_logic;
signal \bfn_14_25_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.running_i\ : std_logic;
signal \current_shift_inst.timer_phase.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.N_192_i\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_2 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_4 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal measured_delay_hc_3 : std_logic;
signal measured_delay_hc_13 : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31\ : std_logic;
signal measured_delay_hc_1 : std_logic;
signal measured_delay_hc_15 : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlt31_0\ : std_logic;
signal measured_delay_hc_8 : std_logic;
signal measured_delay_hc_31 : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_\ : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \current_shift_inst.un4_control_input_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_18\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_30\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_29\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_13\ : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_13 : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_10 : std_logic;
signal \current_shift_inst.N_1742_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_1\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_2\ : std_logic;
signal \current_shift_inst.z_5_2\ : std_logic;
signal \current_shift_inst.z_5_cry_1\ : std_logic;
signal \current_shift_inst.z_5_3\ : std_logic;
signal \current_shift_inst.z_5_cry_2\ : std_logic;
signal \current_shift_inst.z_5_4\ : std_logic;
signal \current_shift_inst.z_5_cry_3\ : std_logic;
signal \current_shift_inst.z_5_5\ : std_logic;
signal \current_shift_inst.z_5_cry_4\ : std_logic;
signal \current_shift_inst.z_5_6\ : std_logic;
signal \current_shift_inst.z_5_cry_5\ : std_logic;
signal \current_shift_inst.z_5_7\ : std_logic;
signal \current_shift_inst.z_5_cry_6\ : std_logic;
signal \current_shift_inst.z_5_8\ : std_logic;
signal \current_shift_inst.z_5_cry_7\ : std_logic;
signal \current_shift_inst.z_5_cry_8\ : std_logic;
signal \current_shift_inst.z_5_9\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \current_shift_inst.z_5_10\ : std_logic;
signal \current_shift_inst.z_5_cry_9\ : std_logic;
signal \current_shift_inst.z_5_11\ : std_logic;
signal \current_shift_inst.z_5_cry_10\ : std_logic;
signal \current_shift_inst.z_5_12\ : std_logic;
signal \current_shift_inst.z_5_cry_11\ : std_logic;
signal \current_shift_inst.z_5_13\ : std_logic;
signal \current_shift_inst.z_5_cry_12\ : std_logic;
signal \current_shift_inst.z_5_14\ : std_logic;
signal \current_shift_inst.z_5_cry_13\ : std_logic;
signal \current_shift_inst.z_5_15\ : std_logic;
signal \current_shift_inst.z_5_cry_14\ : std_logic;
signal \current_shift_inst.z_5_16\ : std_logic;
signal \current_shift_inst.z_5_cry_15\ : std_logic;
signal \current_shift_inst.z_5_cry_16\ : std_logic;
signal \current_shift_inst.z_5_17\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \current_shift_inst.z_5_18\ : std_logic;
signal \current_shift_inst.z_5_cry_17\ : std_logic;
signal \current_shift_inst.z_5_19\ : std_logic;
signal \current_shift_inst.z_5_cry_18\ : std_logic;
signal \current_shift_inst.z_5_20\ : std_logic;
signal \current_shift_inst.z_5_cry_19\ : std_logic;
signal \current_shift_inst.z_5_21\ : std_logic;
signal \current_shift_inst.z_5_cry_20\ : std_logic;
signal \current_shift_inst.z_5_22\ : std_logic;
signal \current_shift_inst.z_5_cry_21\ : std_logic;
signal \current_shift_inst.z_5_23\ : std_logic;
signal \current_shift_inst.z_5_cry_22\ : std_logic;
signal \current_shift_inst.z_5_24\ : std_logic;
signal \current_shift_inst.z_5_cry_23\ : std_logic;
signal \current_shift_inst.z_5_cry_24\ : std_logic;
signal \current_shift_inst.z_5_25\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \current_shift_inst.z_5_26\ : std_logic;
signal \current_shift_inst.z_5_cry_25\ : std_logic;
signal \current_shift_inst.z_5_27\ : std_logic;
signal \current_shift_inst.z_5_cry_26\ : std_logic;
signal \current_shift_inst.z_5_28\ : std_logic;
signal \current_shift_inst.z_5_cry_27\ : std_logic;
signal \current_shift_inst.z_5_29\ : std_logic;
signal \current_shift_inst.z_5_cry_28\ : std_logic;
signal \current_shift_inst.z_5_30\ : std_logic;
signal \current_shift_inst.z_5_cry_29\ : std_logic;
signal \current_shift_inst.z_5_cry_30\ : std_logic;
signal \current_shift_inst.z_5_cry_30_THRU_CO\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\ : std_logic;
signal measured_delay_tr_3 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_20_li\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal measured_delay_tr_8 : std_logic;
signal measured_delay_tr_7 : std_logic;
signal measured_delay_tr_6 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\ : std_logic;
signal measured_delay_tr_5 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_16_17_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_187_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal measured_delay_tr_18 : std_logic;
signal measured_delay_tr_17 : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.N_221_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_424_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_3\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_4\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_5\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_6\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_7\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_8\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_9\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_10\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_11\ : std_logic;
signal \bfn_16_23_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_12\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_13\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_14\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_15\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_16\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_17\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_18\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_19\ : std_logic;
signal \bfn_16_24_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_20\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_21\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_22\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_23\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_24\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_25\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_26\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_27\ : std_logic;
signal \bfn_16_25_0_\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_28\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_29\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_phase.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_30\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_phase_31\ : std_logic;
signal \current_shift_inst.timer_phase.N_188_i_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19\ : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.N_214_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_17_14_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_191_i\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_14\ : std_logic;
signal \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_axb_24\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_390_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_379\ : std_logic;
signal \delay_measurement_inst.N_280_i\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\ : std_logic;
signal \delay_measurement_inst.N_409_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_339_i\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_18_8_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_18_9_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \bfn_18_10_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal s4_phy_c : std_logic;
signal \phase_controller_slave.stateZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.N_213\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal shift_flag_start : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal measured_delay_tr_4 : std_logic;
signal \delay_measurement_inst.N_425\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\ : std_logic;
signal measured_delay_tr_2 : std_logic;
signal \delay_measurement_inst.N_280_i_0\ : std_logic;
signal \delay_measurement_inst.N_286_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_415\ : std_logic;
signal \delay_measurement_inst.N_373\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_18_23_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_18_24_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \bfn_18_25_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_18_26_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.N_211\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_338_i\ : std_logic;
signal red_c_g : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\ <= '0'&\N__18516\&\N__18544\&\N__18517\&\N__18545\&\N__18518\&\N__18174\&\N__18582\&\N__18423\&\N__19705\&\N__18152\&\N__18239\&\N__18319\&\N__18330\&\N__18277\&\N__18288\;
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__43341\&\N__43338\&'0'&'0'&'0'&\N__43336\&\N__43340\&\N__43337\&\N__43339\;
    \pwm_generator_inst.un2_threshold_acc_1_25\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_acc_1_24\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_acc_1_23\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_acc_1_22\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_acc_1_21\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_acc_1_20\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_acc_1_19\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_acc_1_18\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_acc_1_17\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_acc_1_16\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_1_15\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold_acc\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__18552\&\N__18486\&\N__18550\&\N__18485\&\N__18551\&\N__18484\&\N__18553\&\N__18481\&\N__18546\&\N__18480\&\N__18547\&\N__18482\&\N__18548\&\N__18483\&\N__18549\;
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__43500\&\N__43497\&'0'&'0'&'0'&\N__43495\&\N__43499\&\N__43496\&\N__43498\;
    \pwm_generator_inst.un2_threshold_acc_2_1_16\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_acc_2_1_15\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_acc_2_14\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_acc_2_13\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_acc_2_12\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_acc_2_11\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_acc_2_10\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_acc_2_9\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_acc_2_8\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_acc_2_7\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_acc_2_6\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_acc_2_5\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_acc_2_4\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_acc_2_3\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_acc_2_2\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_acc_2_1\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_acc_2_0\ <= \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__20536\,
            RESETB => \N__31431\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43473\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43335\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__43501\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__43494\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__49352\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49354\,
            DIN => \N__49353\,
            DOUT => \N__49352\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49354\,
            PADOUT => \N__49353\,
            PADIN => \N__49352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49343\,
            DIN => \N__49342\,
            DOUT => \N__49341\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49343\,
            PADOUT => \N__49342\,
            PADIN => \N__49341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49334\,
            DIN => \N__49333\,
            DOUT => \N__49332\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49334\,
            PADOUT => \N__49333\,
            PADIN => \N__49332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49325\,
            DIN => \N__49324\,
            DOUT => \N__49323\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49325\,
            PADOUT => \N__49324\,
            PADIN => \N__49323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24697\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49316\,
            DIN => \N__49315\,
            DOUT => \N__49314\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49316\,
            PADOUT => \N__49315\,
            PADIN => \N__49314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49307\,
            DIN => \N__49306\,
            DOUT => \N__49305\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49307\,
            PADOUT => \N__49306\,
            PADIN => \N__49305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49298\,
            DIN => \N__49297\,
            DOUT => \N__49296\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49298\,
            PADOUT => \N__49297\,
            PADIN => \N__49296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49289\,
            DIN => \N__49288\,
            DOUT => \N__49287\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49289\,
            PADOUT => \N__49288\,
            PADIN => \N__49287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49280\,
            DIN => \N__49279\,
            DOUT => \N__49278\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49280\,
            PADOUT => \N__49279\,
            PADIN => \N__49278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49271\,
            DIN => \N__49270\,
            DOUT => \N__49269\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49271\,
            PADOUT => \N__49270\,
            PADIN => \N__49269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30046\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49262\,
            DIN => \N__49261\,
            DOUT => \N__49260\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49262\,
            PADOUT => \N__49261\,
            PADIN => \N__49260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__44785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49253\,
            DIN => \N__49252\,
            DOUT => \N__49251\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__49253\,
            PADOUT => \N__49252\,
            PADIN => \N__49251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__49244\,
            DIN => \N__49243\,
            DOUT => \N__49242\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__49244\,
            PADOUT => \N__49243\,
            PADIN => \N__49242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__45691\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11881\ : InMux
    port map (
            O => \N__49225\,
            I => \N__49221\
        );

    \I__11880\ : InMux
    port map (
            O => \N__49224\,
            I => \N__49218\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__49221\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__11878\ : LocalMux
    port map (
            O => \N__49218\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__11877\ : CascadeMux
    port map (
            O => \N__49213\,
            I => \N__49208\
        );

    \I__11876\ : CascadeMux
    port map (
            O => \N__49212\,
            I => \N__49205\
        );

    \I__11875\ : InMux
    port map (
            O => \N__49211\,
            I => \N__49202\
        );

    \I__11874\ : InMux
    port map (
            O => \N__49208\,
            I => \N__49197\
        );

    \I__11873\ : InMux
    port map (
            O => \N__49205\,
            I => \N__49197\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__49202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__49197\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__11870\ : InMux
    port map (
            O => \N__49192\,
            I => \N__49189\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__49189\,
            I => \N__49186\
        );

    \I__11868\ : Span4Mux_v
    port map (
            O => \N__49186\,
            I => \N__49183\
        );

    \I__11867\ : Odrv4
    port map (
            O => \N__49183\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__11866\ : InMux
    port map (
            O => \N__49180\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__11865\ : InMux
    port map (
            O => \N__49177\,
            I => \N__49173\
        );

    \I__11864\ : InMux
    port map (
            O => \N__49176\,
            I => \N__49170\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__49173\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__49170\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__11861\ : CascadeMux
    port map (
            O => \N__49165\,
            I => \N__49160\
        );

    \I__11860\ : CascadeMux
    port map (
            O => \N__49164\,
            I => \N__49157\
        );

    \I__11859\ : InMux
    port map (
            O => \N__49163\,
            I => \N__49154\
        );

    \I__11858\ : InMux
    port map (
            O => \N__49160\,
            I => \N__49149\
        );

    \I__11857\ : InMux
    port map (
            O => \N__49157\,
            I => \N__49149\
        );

    \I__11856\ : LocalMux
    port map (
            O => \N__49154\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__49149\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__11854\ : InMux
    port map (
            O => \N__49144\,
            I => \N__49141\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__49141\,
            I => \N__49138\
        );

    \I__11852\ : Span4Mux_v
    port map (
            O => \N__49138\,
            I => \N__49135\
        );

    \I__11851\ : Odrv4
    port map (
            O => \N__49135\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__11850\ : InMux
    port map (
            O => \N__49132\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__11849\ : InMux
    port map (
            O => \N__49129\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__11848\ : InMux
    port map (
            O => \N__49126\,
            I => \N__49121\
        );

    \I__11847\ : InMux
    port map (
            O => \N__49125\,
            I => \N__49116\
        );

    \I__11846\ : InMux
    port map (
            O => \N__49124\,
            I => \N__49116\
        );

    \I__11845\ : LocalMux
    port map (
            O => \N__49121\,
            I => \N__49111\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__49116\,
            I => \N__49108\
        );

    \I__11843\ : InMux
    port map (
            O => \N__49115\,
            I => \N__49105\
        );

    \I__11842\ : CascadeMux
    port map (
            O => \N__49114\,
            I => \N__49096\
        );

    \I__11841\ : Span4Mux_h
    port map (
            O => \N__49111\,
            I => \N__49088\
        );

    \I__11840\ : Span4Mux_h
    port map (
            O => \N__49108\,
            I => \N__49088\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__49105\,
            I => \N__49088\
        );

    \I__11838\ : InMux
    port map (
            O => \N__49104\,
            I => \N__49077\
        );

    \I__11837\ : InMux
    port map (
            O => \N__49103\,
            I => \N__49077\
        );

    \I__11836\ : InMux
    port map (
            O => \N__49102\,
            I => \N__49077\
        );

    \I__11835\ : InMux
    port map (
            O => \N__49101\,
            I => \N__49077\
        );

    \I__11834\ : InMux
    port map (
            O => \N__49100\,
            I => \N__49077\
        );

    \I__11833\ : InMux
    port map (
            O => \N__49099\,
            I => \N__49072\
        );

    \I__11832\ : InMux
    port map (
            O => \N__49096\,
            I => \N__49072\
        );

    \I__11831\ : InMux
    port map (
            O => \N__49095\,
            I => \N__49069\
        );

    \I__11830\ : Span4Mux_v
    port map (
            O => \N__49088\,
            I => \N__49066\
        );

    \I__11829\ : LocalMux
    port map (
            O => \N__49077\,
            I => \N__49063\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__49072\,
            I => \N__49058\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__49069\,
            I => \N__49058\
        );

    \I__11826\ : Span4Mux_h
    port map (
            O => \N__49066\,
            I => \N__49053\
        );

    \I__11825\ : Span4Mux_v
    port map (
            O => \N__49063\,
            I => \N__49053\
        );

    \I__11824\ : Span4Mux_v
    port map (
            O => \N__49058\,
            I => \N__49050\
        );

    \I__11823\ : Span4Mux_v
    port map (
            O => \N__49053\,
            I => \N__49047\
        );

    \I__11822\ : Span4Mux_h
    port map (
            O => \N__49050\,
            I => \N__49044\
        );

    \I__11821\ : Odrv4
    port map (
            O => \N__49047\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11820\ : Odrv4
    port map (
            O => \N__49044\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__11819\ : CascadeMux
    port map (
            O => \N__49039\,
            I => \N__49036\
        );

    \I__11818\ : InMux
    port map (
            O => \N__49036\,
            I => \N__49026\
        );

    \I__11817\ : InMux
    port map (
            O => \N__49035\,
            I => \N__49026\
        );

    \I__11816\ : InMux
    port map (
            O => \N__49034\,
            I => \N__49026\
        );

    \I__11815\ : InMux
    port map (
            O => \N__49033\,
            I => \N__49023\
        );

    \I__11814\ : LocalMux
    port map (
            O => \N__49026\,
            I => \N__49018\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__49023\,
            I => \N__49018\
        );

    \I__11812\ : Odrv4
    port map (
            O => \N__49018\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__11811\ : InMux
    port map (
            O => \N__49015\,
            I => \N__49010\
        );

    \I__11810\ : InMux
    port map (
            O => \N__49014\,
            I => \N__49005\
        );

    \I__11809\ : InMux
    port map (
            O => \N__49013\,
            I => \N__49005\
        );

    \I__11808\ : LocalMux
    port map (
            O => \N__49010\,
            I => \N__49002\
        );

    \I__11807\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48999\
        );

    \I__11806\ : Span4Mux_v
    port map (
            O => \N__49002\,
            I => \N__48996\
        );

    \I__11805\ : Span4Mux_v
    port map (
            O => \N__48999\,
            I => \N__48993\
        );

    \I__11804\ : Span4Mux_h
    port map (
            O => \N__48996\,
            I => \N__48990\
        );

    \I__11803\ : Odrv4
    port map (
            O => \N__48993\,
            I => \il_min_comp2_D2\
        );

    \I__11802\ : Odrv4
    port map (
            O => \N__48990\,
            I => \il_min_comp2_D2\
        );

    \I__11801\ : InMux
    port map (
            O => \N__48985\,
            I => \N__48982\
        );

    \I__11800\ : LocalMux
    port map (
            O => \N__48982\,
            I => \N__48979\
        );

    \I__11799\ : Span4Mux_h
    port map (
            O => \N__48979\,
            I => \N__48976\
        );

    \I__11798\ : Odrv4
    port map (
            O => \N__48976\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__11797\ : InMux
    port map (
            O => \N__48973\,
            I => \N__48968\
        );

    \I__11796\ : InMux
    port map (
            O => \N__48972\,
            I => \N__48965\
        );

    \I__11795\ : InMux
    port map (
            O => \N__48971\,
            I => \N__48962\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__48968\,
            I => \N__48959\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__48965\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__48962\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__11791\ : Odrv4
    port map (
            O => \N__48959\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__11790\ : InMux
    port map (
            O => \N__48952\,
            I => \N__48949\
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__48949\,
            I => \N__48945\
        );

    \I__11788\ : InMux
    port map (
            O => \N__48948\,
            I => \N__48942\
        );

    \I__11787\ : Span4Mux_h
    port map (
            O => \N__48945\,
            I => \N__48939\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__48942\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__11785\ : Odrv4
    port map (
            O => \N__48939\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__11784\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48928\
        );

    \I__11783\ : InMux
    port map (
            O => \N__48933\,
            I => \N__48928\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__48928\,
            I => \N__48925\
        );

    \I__11781\ : Odrv4
    port map (
            O => \N__48925\,
            I => \phase_controller_slave.N_211\
        );

    \I__11780\ : InMux
    port map (
            O => \N__48922\,
            I => \N__48919\
        );

    \I__11779\ : LocalMux
    port map (
            O => \N__48919\,
            I => \N__48916\
        );

    \I__11778\ : Span4Mux_v
    port map (
            O => \N__48916\,
            I => \N__48913\
        );

    \I__11777\ : Span4Mux_h
    port map (
            O => \N__48913\,
            I => \N__48908\
        );

    \I__11776\ : InMux
    port map (
            O => \N__48912\,
            I => \N__48905\
        );

    \I__11775\ : InMux
    port map (
            O => \N__48911\,
            I => \N__48902\
        );

    \I__11774\ : Odrv4
    port map (
            O => \N__48908\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11773\ : LocalMux
    port map (
            O => \N__48905\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__48902\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__11771\ : InMux
    port map (
            O => \N__48895\,
            I => \N__48891\
        );

    \I__11770\ : InMux
    port map (
            O => \N__48894\,
            I => \N__48888\
        );

    \I__11769\ : LocalMux
    port map (
            O => \N__48891\,
            I => \N__48885\
        );

    \I__11768\ : LocalMux
    port map (
            O => \N__48888\,
            I => \N__48882\
        );

    \I__11767\ : Span4Mux_h
    port map (
            O => \N__48885\,
            I => \N__48879\
        );

    \I__11766\ : Odrv12
    port map (
            O => \N__48882\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__11765\ : Odrv4
    port map (
            O => \N__48879\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__11764\ : ClkMux
    port map (
            O => \N__48874\,
            I => \N__48349\
        );

    \I__11763\ : ClkMux
    port map (
            O => \N__48873\,
            I => \N__48349\
        );

    \I__11762\ : ClkMux
    port map (
            O => \N__48872\,
            I => \N__48349\
        );

    \I__11761\ : ClkMux
    port map (
            O => \N__48871\,
            I => \N__48349\
        );

    \I__11760\ : ClkMux
    port map (
            O => \N__48870\,
            I => \N__48349\
        );

    \I__11759\ : ClkMux
    port map (
            O => \N__48869\,
            I => \N__48349\
        );

    \I__11758\ : ClkMux
    port map (
            O => \N__48868\,
            I => \N__48349\
        );

    \I__11757\ : ClkMux
    port map (
            O => \N__48867\,
            I => \N__48349\
        );

    \I__11756\ : ClkMux
    port map (
            O => \N__48866\,
            I => \N__48349\
        );

    \I__11755\ : ClkMux
    port map (
            O => \N__48865\,
            I => \N__48349\
        );

    \I__11754\ : ClkMux
    port map (
            O => \N__48864\,
            I => \N__48349\
        );

    \I__11753\ : ClkMux
    port map (
            O => \N__48863\,
            I => \N__48349\
        );

    \I__11752\ : ClkMux
    port map (
            O => \N__48862\,
            I => \N__48349\
        );

    \I__11751\ : ClkMux
    port map (
            O => \N__48861\,
            I => \N__48349\
        );

    \I__11750\ : ClkMux
    port map (
            O => \N__48860\,
            I => \N__48349\
        );

    \I__11749\ : ClkMux
    port map (
            O => \N__48859\,
            I => \N__48349\
        );

    \I__11748\ : ClkMux
    port map (
            O => \N__48858\,
            I => \N__48349\
        );

    \I__11747\ : ClkMux
    port map (
            O => \N__48857\,
            I => \N__48349\
        );

    \I__11746\ : ClkMux
    port map (
            O => \N__48856\,
            I => \N__48349\
        );

    \I__11745\ : ClkMux
    port map (
            O => \N__48855\,
            I => \N__48349\
        );

    \I__11744\ : ClkMux
    port map (
            O => \N__48854\,
            I => \N__48349\
        );

    \I__11743\ : ClkMux
    port map (
            O => \N__48853\,
            I => \N__48349\
        );

    \I__11742\ : ClkMux
    port map (
            O => \N__48852\,
            I => \N__48349\
        );

    \I__11741\ : ClkMux
    port map (
            O => \N__48851\,
            I => \N__48349\
        );

    \I__11740\ : ClkMux
    port map (
            O => \N__48850\,
            I => \N__48349\
        );

    \I__11739\ : ClkMux
    port map (
            O => \N__48849\,
            I => \N__48349\
        );

    \I__11738\ : ClkMux
    port map (
            O => \N__48848\,
            I => \N__48349\
        );

    \I__11737\ : ClkMux
    port map (
            O => \N__48847\,
            I => \N__48349\
        );

    \I__11736\ : ClkMux
    port map (
            O => \N__48846\,
            I => \N__48349\
        );

    \I__11735\ : ClkMux
    port map (
            O => \N__48845\,
            I => \N__48349\
        );

    \I__11734\ : ClkMux
    port map (
            O => \N__48844\,
            I => \N__48349\
        );

    \I__11733\ : ClkMux
    port map (
            O => \N__48843\,
            I => \N__48349\
        );

    \I__11732\ : ClkMux
    port map (
            O => \N__48842\,
            I => \N__48349\
        );

    \I__11731\ : ClkMux
    port map (
            O => \N__48841\,
            I => \N__48349\
        );

    \I__11730\ : ClkMux
    port map (
            O => \N__48840\,
            I => \N__48349\
        );

    \I__11729\ : ClkMux
    port map (
            O => \N__48839\,
            I => \N__48349\
        );

    \I__11728\ : ClkMux
    port map (
            O => \N__48838\,
            I => \N__48349\
        );

    \I__11727\ : ClkMux
    port map (
            O => \N__48837\,
            I => \N__48349\
        );

    \I__11726\ : ClkMux
    port map (
            O => \N__48836\,
            I => \N__48349\
        );

    \I__11725\ : ClkMux
    port map (
            O => \N__48835\,
            I => \N__48349\
        );

    \I__11724\ : ClkMux
    port map (
            O => \N__48834\,
            I => \N__48349\
        );

    \I__11723\ : ClkMux
    port map (
            O => \N__48833\,
            I => \N__48349\
        );

    \I__11722\ : ClkMux
    port map (
            O => \N__48832\,
            I => \N__48349\
        );

    \I__11721\ : ClkMux
    port map (
            O => \N__48831\,
            I => \N__48349\
        );

    \I__11720\ : ClkMux
    port map (
            O => \N__48830\,
            I => \N__48349\
        );

    \I__11719\ : ClkMux
    port map (
            O => \N__48829\,
            I => \N__48349\
        );

    \I__11718\ : ClkMux
    port map (
            O => \N__48828\,
            I => \N__48349\
        );

    \I__11717\ : ClkMux
    port map (
            O => \N__48827\,
            I => \N__48349\
        );

    \I__11716\ : ClkMux
    port map (
            O => \N__48826\,
            I => \N__48349\
        );

    \I__11715\ : ClkMux
    port map (
            O => \N__48825\,
            I => \N__48349\
        );

    \I__11714\ : ClkMux
    port map (
            O => \N__48824\,
            I => \N__48349\
        );

    \I__11713\ : ClkMux
    port map (
            O => \N__48823\,
            I => \N__48349\
        );

    \I__11712\ : ClkMux
    port map (
            O => \N__48822\,
            I => \N__48349\
        );

    \I__11711\ : ClkMux
    port map (
            O => \N__48821\,
            I => \N__48349\
        );

    \I__11710\ : ClkMux
    port map (
            O => \N__48820\,
            I => \N__48349\
        );

    \I__11709\ : ClkMux
    port map (
            O => \N__48819\,
            I => \N__48349\
        );

    \I__11708\ : ClkMux
    port map (
            O => \N__48818\,
            I => \N__48349\
        );

    \I__11707\ : ClkMux
    port map (
            O => \N__48817\,
            I => \N__48349\
        );

    \I__11706\ : ClkMux
    port map (
            O => \N__48816\,
            I => \N__48349\
        );

    \I__11705\ : ClkMux
    port map (
            O => \N__48815\,
            I => \N__48349\
        );

    \I__11704\ : ClkMux
    port map (
            O => \N__48814\,
            I => \N__48349\
        );

    \I__11703\ : ClkMux
    port map (
            O => \N__48813\,
            I => \N__48349\
        );

    \I__11702\ : ClkMux
    port map (
            O => \N__48812\,
            I => \N__48349\
        );

    \I__11701\ : ClkMux
    port map (
            O => \N__48811\,
            I => \N__48349\
        );

    \I__11700\ : ClkMux
    port map (
            O => \N__48810\,
            I => \N__48349\
        );

    \I__11699\ : ClkMux
    port map (
            O => \N__48809\,
            I => \N__48349\
        );

    \I__11698\ : ClkMux
    port map (
            O => \N__48808\,
            I => \N__48349\
        );

    \I__11697\ : ClkMux
    port map (
            O => \N__48807\,
            I => \N__48349\
        );

    \I__11696\ : ClkMux
    port map (
            O => \N__48806\,
            I => \N__48349\
        );

    \I__11695\ : ClkMux
    port map (
            O => \N__48805\,
            I => \N__48349\
        );

    \I__11694\ : ClkMux
    port map (
            O => \N__48804\,
            I => \N__48349\
        );

    \I__11693\ : ClkMux
    port map (
            O => \N__48803\,
            I => \N__48349\
        );

    \I__11692\ : ClkMux
    port map (
            O => \N__48802\,
            I => \N__48349\
        );

    \I__11691\ : ClkMux
    port map (
            O => \N__48801\,
            I => \N__48349\
        );

    \I__11690\ : ClkMux
    port map (
            O => \N__48800\,
            I => \N__48349\
        );

    \I__11689\ : ClkMux
    port map (
            O => \N__48799\,
            I => \N__48349\
        );

    \I__11688\ : ClkMux
    port map (
            O => \N__48798\,
            I => \N__48349\
        );

    \I__11687\ : ClkMux
    port map (
            O => \N__48797\,
            I => \N__48349\
        );

    \I__11686\ : ClkMux
    port map (
            O => \N__48796\,
            I => \N__48349\
        );

    \I__11685\ : ClkMux
    port map (
            O => \N__48795\,
            I => \N__48349\
        );

    \I__11684\ : ClkMux
    port map (
            O => \N__48794\,
            I => \N__48349\
        );

    \I__11683\ : ClkMux
    port map (
            O => \N__48793\,
            I => \N__48349\
        );

    \I__11682\ : ClkMux
    port map (
            O => \N__48792\,
            I => \N__48349\
        );

    \I__11681\ : ClkMux
    port map (
            O => \N__48791\,
            I => \N__48349\
        );

    \I__11680\ : ClkMux
    port map (
            O => \N__48790\,
            I => \N__48349\
        );

    \I__11679\ : ClkMux
    port map (
            O => \N__48789\,
            I => \N__48349\
        );

    \I__11678\ : ClkMux
    port map (
            O => \N__48788\,
            I => \N__48349\
        );

    \I__11677\ : ClkMux
    port map (
            O => \N__48787\,
            I => \N__48349\
        );

    \I__11676\ : ClkMux
    port map (
            O => \N__48786\,
            I => \N__48349\
        );

    \I__11675\ : ClkMux
    port map (
            O => \N__48785\,
            I => \N__48349\
        );

    \I__11674\ : ClkMux
    port map (
            O => \N__48784\,
            I => \N__48349\
        );

    \I__11673\ : ClkMux
    port map (
            O => \N__48783\,
            I => \N__48349\
        );

    \I__11672\ : ClkMux
    port map (
            O => \N__48782\,
            I => \N__48349\
        );

    \I__11671\ : ClkMux
    port map (
            O => \N__48781\,
            I => \N__48349\
        );

    \I__11670\ : ClkMux
    port map (
            O => \N__48780\,
            I => \N__48349\
        );

    \I__11669\ : ClkMux
    port map (
            O => \N__48779\,
            I => \N__48349\
        );

    \I__11668\ : ClkMux
    port map (
            O => \N__48778\,
            I => \N__48349\
        );

    \I__11667\ : ClkMux
    port map (
            O => \N__48777\,
            I => \N__48349\
        );

    \I__11666\ : ClkMux
    port map (
            O => \N__48776\,
            I => \N__48349\
        );

    \I__11665\ : ClkMux
    port map (
            O => \N__48775\,
            I => \N__48349\
        );

    \I__11664\ : ClkMux
    port map (
            O => \N__48774\,
            I => \N__48349\
        );

    \I__11663\ : ClkMux
    port map (
            O => \N__48773\,
            I => \N__48349\
        );

    \I__11662\ : ClkMux
    port map (
            O => \N__48772\,
            I => \N__48349\
        );

    \I__11661\ : ClkMux
    port map (
            O => \N__48771\,
            I => \N__48349\
        );

    \I__11660\ : ClkMux
    port map (
            O => \N__48770\,
            I => \N__48349\
        );

    \I__11659\ : ClkMux
    port map (
            O => \N__48769\,
            I => \N__48349\
        );

    \I__11658\ : ClkMux
    port map (
            O => \N__48768\,
            I => \N__48349\
        );

    \I__11657\ : ClkMux
    port map (
            O => \N__48767\,
            I => \N__48349\
        );

    \I__11656\ : ClkMux
    port map (
            O => \N__48766\,
            I => \N__48349\
        );

    \I__11655\ : ClkMux
    port map (
            O => \N__48765\,
            I => \N__48349\
        );

    \I__11654\ : ClkMux
    port map (
            O => \N__48764\,
            I => \N__48349\
        );

    \I__11653\ : ClkMux
    port map (
            O => \N__48763\,
            I => \N__48349\
        );

    \I__11652\ : ClkMux
    port map (
            O => \N__48762\,
            I => \N__48349\
        );

    \I__11651\ : ClkMux
    port map (
            O => \N__48761\,
            I => \N__48349\
        );

    \I__11650\ : ClkMux
    port map (
            O => \N__48760\,
            I => \N__48349\
        );

    \I__11649\ : ClkMux
    port map (
            O => \N__48759\,
            I => \N__48349\
        );

    \I__11648\ : ClkMux
    port map (
            O => \N__48758\,
            I => \N__48349\
        );

    \I__11647\ : ClkMux
    port map (
            O => \N__48757\,
            I => \N__48349\
        );

    \I__11646\ : ClkMux
    port map (
            O => \N__48756\,
            I => \N__48349\
        );

    \I__11645\ : ClkMux
    port map (
            O => \N__48755\,
            I => \N__48349\
        );

    \I__11644\ : ClkMux
    port map (
            O => \N__48754\,
            I => \N__48349\
        );

    \I__11643\ : ClkMux
    port map (
            O => \N__48753\,
            I => \N__48349\
        );

    \I__11642\ : ClkMux
    port map (
            O => \N__48752\,
            I => \N__48349\
        );

    \I__11641\ : ClkMux
    port map (
            O => \N__48751\,
            I => \N__48349\
        );

    \I__11640\ : ClkMux
    port map (
            O => \N__48750\,
            I => \N__48349\
        );

    \I__11639\ : ClkMux
    port map (
            O => \N__48749\,
            I => \N__48349\
        );

    \I__11638\ : ClkMux
    port map (
            O => \N__48748\,
            I => \N__48349\
        );

    \I__11637\ : ClkMux
    port map (
            O => \N__48747\,
            I => \N__48349\
        );

    \I__11636\ : ClkMux
    port map (
            O => \N__48746\,
            I => \N__48349\
        );

    \I__11635\ : ClkMux
    port map (
            O => \N__48745\,
            I => \N__48349\
        );

    \I__11634\ : ClkMux
    port map (
            O => \N__48744\,
            I => \N__48349\
        );

    \I__11633\ : ClkMux
    port map (
            O => \N__48743\,
            I => \N__48349\
        );

    \I__11632\ : ClkMux
    port map (
            O => \N__48742\,
            I => \N__48349\
        );

    \I__11631\ : ClkMux
    port map (
            O => \N__48741\,
            I => \N__48349\
        );

    \I__11630\ : ClkMux
    port map (
            O => \N__48740\,
            I => \N__48349\
        );

    \I__11629\ : ClkMux
    port map (
            O => \N__48739\,
            I => \N__48349\
        );

    \I__11628\ : ClkMux
    port map (
            O => \N__48738\,
            I => \N__48349\
        );

    \I__11627\ : ClkMux
    port map (
            O => \N__48737\,
            I => \N__48349\
        );

    \I__11626\ : ClkMux
    port map (
            O => \N__48736\,
            I => \N__48349\
        );

    \I__11625\ : ClkMux
    port map (
            O => \N__48735\,
            I => \N__48349\
        );

    \I__11624\ : ClkMux
    port map (
            O => \N__48734\,
            I => \N__48349\
        );

    \I__11623\ : ClkMux
    port map (
            O => \N__48733\,
            I => \N__48349\
        );

    \I__11622\ : ClkMux
    port map (
            O => \N__48732\,
            I => \N__48349\
        );

    \I__11621\ : ClkMux
    port map (
            O => \N__48731\,
            I => \N__48349\
        );

    \I__11620\ : ClkMux
    port map (
            O => \N__48730\,
            I => \N__48349\
        );

    \I__11619\ : ClkMux
    port map (
            O => \N__48729\,
            I => \N__48349\
        );

    \I__11618\ : ClkMux
    port map (
            O => \N__48728\,
            I => \N__48349\
        );

    \I__11617\ : ClkMux
    port map (
            O => \N__48727\,
            I => \N__48349\
        );

    \I__11616\ : ClkMux
    port map (
            O => \N__48726\,
            I => \N__48349\
        );

    \I__11615\ : ClkMux
    port map (
            O => \N__48725\,
            I => \N__48349\
        );

    \I__11614\ : ClkMux
    port map (
            O => \N__48724\,
            I => \N__48349\
        );

    \I__11613\ : ClkMux
    port map (
            O => \N__48723\,
            I => \N__48349\
        );

    \I__11612\ : ClkMux
    port map (
            O => \N__48722\,
            I => \N__48349\
        );

    \I__11611\ : ClkMux
    port map (
            O => \N__48721\,
            I => \N__48349\
        );

    \I__11610\ : ClkMux
    port map (
            O => \N__48720\,
            I => \N__48349\
        );

    \I__11609\ : ClkMux
    port map (
            O => \N__48719\,
            I => \N__48349\
        );

    \I__11608\ : ClkMux
    port map (
            O => \N__48718\,
            I => \N__48349\
        );

    \I__11607\ : ClkMux
    port map (
            O => \N__48717\,
            I => \N__48349\
        );

    \I__11606\ : ClkMux
    port map (
            O => \N__48716\,
            I => \N__48349\
        );

    \I__11605\ : ClkMux
    port map (
            O => \N__48715\,
            I => \N__48349\
        );

    \I__11604\ : ClkMux
    port map (
            O => \N__48714\,
            I => \N__48349\
        );

    \I__11603\ : ClkMux
    port map (
            O => \N__48713\,
            I => \N__48349\
        );

    \I__11602\ : ClkMux
    port map (
            O => \N__48712\,
            I => \N__48349\
        );

    \I__11601\ : ClkMux
    port map (
            O => \N__48711\,
            I => \N__48349\
        );

    \I__11600\ : ClkMux
    port map (
            O => \N__48710\,
            I => \N__48349\
        );

    \I__11599\ : ClkMux
    port map (
            O => \N__48709\,
            I => \N__48349\
        );

    \I__11598\ : ClkMux
    port map (
            O => \N__48708\,
            I => \N__48349\
        );

    \I__11597\ : ClkMux
    port map (
            O => \N__48707\,
            I => \N__48349\
        );

    \I__11596\ : ClkMux
    port map (
            O => \N__48706\,
            I => \N__48349\
        );

    \I__11595\ : ClkMux
    port map (
            O => \N__48705\,
            I => \N__48349\
        );

    \I__11594\ : ClkMux
    port map (
            O => \N__48704\,
            I => \N__48349\
        );

    \I__11593\ : ClkMux
    port map (
            O => \N__48703\,
            I => \N__48349\
        );

    \I__11592\ : ClkMux
    port map (
            O => \N__48702\,
            I => \N__48349\
        );

    \I__11591\ : ClkMux
    port map (
            O => \N__48701\,
            I => \N__48349\
        );

    \I__11590\ : ClkMux
    port map (
            O => \N__48700\,
            I => \N__48349\
        );

    \I__11589\ : GlobalMux
    port map (
            O => \N__48349\,
            I => clk_100mhz_0
        );

    \I__11588\ : CEMux
    port map (
            O => \N__48346\,
            I => \N__48340\
        );

    \I__11587\ : CEMux
    port map (
            O => \N__48345\,
            I => \N__48335\
        );

    \I__11586\ : CEMux
    port map (
            O => \N__48344\,
            I => \N__48332\
        );

    \I__11585\ : CEMux
    port map (
            O => \N__48343\,
            I => \N__48329\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__48340\,
            I => \N__48326\
        );

    \I__11583\ : CEMux
    port map (
            O => \N__48339\,
            I => \N__48323\
        );

    \I__11582\ : CEMux
    port map (
            O => \N__48338\,
            I => \N__48320\
        );

    \I__11581\ : LocalMux
    port map (
            O => \N__48335\,
            I => \N__48317\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__48332\,
            I => \N__48312\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__48329\,
            I => \N__48312\
        );

    \I__11578\ : Span4Mux_h
    port map (
            O => \N__48326\,
            I => \N__48309\
        );

    \I__11577\ : LocalMux
    port map (
            O => \N__48323\,
            I => \N__48306\
        );

    \I__11576\ : LocalMux
    port map (
            O => \N__48320\,
            I => \N__48303\
        );

    \I__11575\ : Span12Mux_s8_h
    port map (
            O => \N__48317\,
            I => \N__48300\
        );

    \I__11574\ : Span4Mux_v
    port map (
            O => \N__48312\,
            I => \N__48297\
        );

    \I__11573\ : Span4Mux_v
    port map (
            O => \N__48309\,
            I => \N__48292\
        );

    \I__11572\ : Span4Mux_v
    port map (
            O => \N__48306\,
            I => \N__48292\
        );

    \I__11571\ : Span4Mux_h
    port map (
            O => \N__48303\,
            I => \N__48289\
        );

    \I__11570\ : Odrv12
    port map (
            O => \N__48300\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__11569\ : Odrv4
    port map (
            O => \N__48297\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__11568\ : Odrv4
    port map (
            O => \N__48292\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__11567\ : Odrv4
    port map (
            O => \N__48289\,
            I => \delay_measurement_inst.delay_tr_timer.N_338_i\
        );

    \I__11566\ : CascadeMux
    port map (
            O => \N__48280\,
            I => \N__48272\
        );

    \I__11565\ : InMux
    port map (
            O => \N__48279\,
            I => \N__48269\
        );

    \I__11564\ : InMux
    port map (
            O => \N__48278\,
            I => \N__48266\
        );

    \I__11563\ : InMux
    port map (
            O => \N__48277\,
            I => \N__48263\
        );

    \I__11562\ : InMux
    port map (
            O => \N__48276\,
            I => \N__48260\
        );

    \I__11561\ : InMux
    port map (
            O => \N__48275\,
            I => \N__48257\
        );

    \I__11560\ : InMux
    port map (
            O => \N__48272\,
            I => \N__48254\
        );

    \I__11559\ : LocalMux
    port map (
            O => \N__48269\,
            I => \N__48251\
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__48266\,
            I => \N__48248\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__48263\,
            I => \N__48245\
        );

    \I__11556\ : LocalMux
    port map (
            O => \N__48260\,
            I => \N__48242\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__48257\,
            I => \N__48167\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__48254\,
            I => \N__48114\
        );

    \I__11553\ : Glb2LocalMux
    port map (
            O => \N__48251\,
            I => \N__47779\
        );

    \I__11552\ : Glb2LocalMux
    port map (
            O => \N__48248\,
            I => \N__47779\
        );

    \I__11551\ : Glb2LocalMux
    port map (
            O => \N__48245\,
            I => \N__47779\
        );

    \I__11550\ : Glb2LocalMux
    port map (
            O => \N__48242\,
            I => \N__47779\
        );

    \I__11549\ : SRMux
    port map (
            O => \N__48241\,
            I => \N__47779\
        );

    \I__11548\ : SRMux
    port map (
            O => \N__48240\,
            I => \N__47779\
        );

    \I__11547\ : SRMux
    port map (
            O => \N__48239\,
            I => \N__47779\
        );

    \I__11546\ : SRMux
    port map (
            O => \N__48238\,
            I => \N__47779\
        );

    \I__11545\ : SRMux
    port map (
            O => \N__48237\,
            I => \N__47779\
        );

    \I__11544\ : SRMux
    port map (
            O => \N__48236\,
            I => \N__47779\
        );

    \I__11543\ : SRMux
    port map (
            O => \N__48235\,
            I => \N__47779\
        );

    \I__11542\ : SRMux
    port map (
            O => \N__48234\,
            I => \N__47779\
        );

    \I__11541\ : SRMux
    port map (
            O => \N__48233\,
            I => \N__47779\
        );

    \I__11540\ : SRMux
    port map (
            O => \N__48232\,
            I => \N__47779\
        );

    \I__11539\ : SRMux
    port map (
            O => \N__48231\,
            I => \N__47779\
        );

    \I__11538\ : SRMux
    port map (
            O => \N__48230\,
            I => \N__47779\
        );

    \I__11537\ : SRMux
    port map (
            O => \N__48229\,
            I => \N__47779\
        );

    \I__11536\ : SRMux
    port map (
            O => \N__48228\,
            I => \N__47779\
        );

    \I__11535\ : SRMux
    port map (
            O => \N__48227\,
            I => \N__47779\
        );

    \I__11534\ : SRMux
    port map (
            O => \N__48226\,
            I => \N__47779\
        );

    \I__11533\ : SRMux
    port map (
            O => \N__48225\,
            I => \N__47779\
        );

    \I__11532\ : SRMux
    port map (
            O => \N__48224\,
            I => \N__47779\
        );

    \I__11531\ : SRMux
    port map (
            O => \N__48223\,
            I => \N__47779\
        );

    \I__11530\ : SRMux
    port map (
            O => \N__48222\,
            I => \N__47779\
        );

    \I__11529\ : SRMux
    port map (
            O => \N__48221\,
            I => \N__47779\
        );

    \I__11528\ : SRMux
    port map (
            O => \N__48220\,
            I => \N__47779\
        );

    \I__11527\ : SRMux
    port map (
            O => \N__48219\,
            I => \N__47779\
        );

    \I__11526\ : SRMux
    port map (
            O => \N__48218\,
            I => \N__47779\
        );

    \I__11525\ : SRMux
    port map (
            O => \N__48217\,
            I => \N__47779\
        );

    \I__11524\ : SRMux
    port map (
            O => \N__48216\,
            I => \N__47779\
        );

    \I__11523\ : SRMux
    port map (
            O => \N__48215\,
            I => \N__47779\
        );

    \I__11522\ : SRMux
    port map (
            O => \N__48214\,
            I => \N__47779\
        );

    \I__11521\ : SRMux
    port map (
            O => \N__48213\,
            I => \N__47779\
        );

    \I__11520\ : SRMux
    port map (
            O => \N__48212\,
            I => \N__47779\
        );

    \I__11519\ : SRMux
    port map (
            O => \N__48211\,
            I => \N__47779\
        );

    \I__11518\ : SRMux
    port map (
            O => \N__48210\,
            I => \N__47779\
        );

    \I__11517\ : SRMux
    port map (
            O => \N__48209\,
            I => \N__47779\
        );

    \I__11516\ : SRMux
    port map (
            O => \N__48208\,
            I => \N__47779\
        );

    \I__11515\ : SRMux
    port map (
            O => \N__48207\,
            I => \N__47779\
        );

    \I__11514\ : SRMux
    port map (
            O => \N__48206\,
            I => \N__47779\
        );

    \I__11513\ : SRMux
    port map (
            O => \N__48205\,
            I => \N__47779\
        );

    \I__11512\ : SRMux
    port map (
            O => \N__48204\,
            I => \N__47779\
        );

    \I__11511\ : SRMux
    port map (
            O => \N__48203\,
            I => \N__47779\
        );

    \I__11510\ : SRMux
    port map (
            O => \N__48202\,
            I => \N__47779\
        );

    \I__11509\ : SRMux
    port map (
            O => \N__48201\,
            I => \N__47779\
        );

    \I__11508\ : SRMux
    port map (
            O => \N__48200\,
            I => \N__47779\
        );

    \I__11507\ : SRMux
    port map (
            O => \N__48199\,
            I => \N__47779\
        );

    \I__11506\ : SRMux
    port map (
            O => \N__48198\,
            I => \N__47779\
        );

    \I__11505\ : SRMux
    port map (
            O => \N__48197\,
            I => \N__47779\
        );

    \I__11504\ : SRMux
    port map (
            O => \N__48196\,
            I => \N__47779\
        );

    \I__11503\ : SRMux
    port map (
            O => \N__48195\,
            I => \N__47779\
        );

    \I__11502\ : SRMux
    port map (
            O => \N__48194\,
            I => \N__47779\
        );

    \I__11501\ : SRMux
    port map (
            O => \N__48193\,
            I => \N__47779\
        );

    \I__11500\ : SRMux
    port map (
            O => \N__48192\,
            I => \N__47779\
        );

    \I__11499\ : SRMux
    port map (
            O => \N__48191\,
            I => \N__47779\
        );

    \I__11498\ : SRMux
    port map (
            O => \N__48190\,
            I => \N__47779\
        );

    \I__11497\ : SRMux
    port map (
            O => \N__48189\,
            I => \N__47779\
        );

    \I__11496\ : SRMux
    port map (
            O => \N__48188\,
            I => \N__47779\
        );

    \I__11495\ : SRMux
    port map (
            O => \N__48187\,
            I => \N__47779\
        );

    \I__11494\ : SRMux
    port map (
            O => \N__48186\,
            I => \N__47779\
        );

    \I__11493\ : SRMux
    port map (
            O => \N__48185\,
            I => \N__47779\
        );

    \I__11492\ : SRMux
    port map (
            O => \N__48184\,
            I => \N__47779\
        );

    \I__11491\ : SRMux
    port map (
            O => \N__48183\,
            I => \N__47779\
        );

    \I__11490\ : SRMux
    port map (
            O => \N__48182\,
            I => \N__47779\
        );

    \I__11489\ : SRMux
    port map (
            O => \N__48181\,
            I => \N__47779\
        );

    \I__11488\ : SRMux
    port map (
            O => \N__48180\,
            I => \N__47779\
        );

    \I__11487\ : SRMux
    port map (
            O => \N__48179\,
            I => \N__47779\
        );

    \I__11486\ : SRMux
    port map (
            O => \N__48178\,
            I => \N__47779\
        );

    \I__11485\ : SRMux
    port map (
            O => \N__48177\,
            I => \N__47779\
        );

    \I__11484\ : SRMux
    port map (
            O => \N__48176\,
            I => \N__47779\
        );

    \I__11483\ : SRMux
    port map (
            O => \N__48175\,
            I => \N__47779\
        );

    \I__11482\ : SRMux
    port map (
            O => \N__48174\,
            I => \N__47779\
        );

    \I__11481\ : SRMux
    port map (
            O => \N__48173\,
            I => \N__47779\
        );

    \I__11480\ : SRMux
    port map (
            O => \N__48172\,
            I => \N__47779\
        );

    \I__11479\ : SRMux
    port map (
            O => \N__48171\,
            I => \N__47779\
        );

    \I__11478\ : SRMux
    port map (
            O => \N__48170\,
            I => \N__47779\
        );

    \I__11477\ : Glb2LocalMux
    port map (
            O => \N__48167\,
            I => \N__47779\
        );

    \I__11476\ : SRMux
    port map (
            O => \N__48166\,
            I => \N__47779\
        );

    \I__11475\ : SRMux
    port map (
            O => \N__48165\,
            I => \N__47779\
        );

    \I__11474\ : SRMux
    port map (
            O => \N__48164\,
            I => \N__47779\
        );

    \I__11473\ : SRMux
    port map (
            O => \N__48163\,
            I => \N__47779\
        );

    \I__11472\ : SRMux
    port map (
            O => \N__48162\,
            I => \N__47779\
        );

    \I__11471\ : SRMux
    port map (
            O => \N__48161\,
            I => \N__47779\
        );

    \I__11470\ : SRMux
    port map (
            O => \N__48160\,
            I => \N__47779\
        );

    \I__11469\ : SRMux
    port map (
            O => \N__48159\,
            I => \N__47779\
        );

    \I__11468\ : SRMux
    port map (
            O => \N__48158\,
            I => \N__47779\
        );

    \I__11467\ : SRMux
    port map (
            O => \N__48157\,
            I => \N__47779\
        );

    \I__11466\ : SRMux
    port map (
            O => \N__48156\,
            I => \N__47779\
        );

    \I__11465\ : SRMux
    port map (
            O => \N__48155\,
            I => \N__47779\
        );

    \I__11464\ : SRMux
    port map (
            O => \N__48154\,
            I => \N__47779\
        );

    \I__11463\ : SRMux
    port map (
            O => \N__48153\,
            I => \N__47779\
        );

    \I__11462\ : SRMux
    port map (
            O => \N__48152\,
            I => \N__47779\
        );

    \I__11461\ : SRMux
    port map (
            O => \N__48151\,
            I => \N__47779\
        );

    \I__11460\ : SRMux
    port map (
            O => \N__48150\,
            I => \N__47779\
        );

    \I__11459\ : SRMux
    port map (
            O => \N__48149\,
            I => \N__47779\
        );

    \I__11458\ : SRMux
    port map (
            O => \N__48148\,
            I => \N__47779\
        );

    \I__11457\ : SRMux
    port map (
            O => \N__48147\,
            I => \N__47779\
        );

    \I__11456\ : SRMux
    port map (
            O => \N__48146\,
            I => \N__47779\
        );

    \I__11455\ : SRMux
    port map (
            O => \N__48145\,
            I => \N__47779\
        );

    \I__11454\ : SRMux
    port map (
            O => \N__48144\,
            I => \N__47779\
        );

    \I__11453\ : SRMux
    port map (
            O => \N__48143\,
            I => \N__47779\
        );

    \I__11452\ : SRMux
    port map (
            O => \N__48142\,
            I => \N__47779\
        );

    \I__11451\ : SRMux
    port map (
            O => \N__48141\,
            I => \N__47779\
        );

    \I__11450\ : SRMux
    port map (
            O => \N__48140\,
            I => \N__47779\
        );

    \I__11449\ : SRMux
    port map (
            O => \N__48139\,
            I => \N__47779\
        );

    \I__11448\ : SRMux
    port map (
            O => \N__48138\,
            I => \N__47779\
        );

    \I__11447\ : SRMux
    port map (
            O => \N__48137\,
            I => \N__47779\
        );

    \I__11446\ : SRMux
    port map (
            O => \N__48136\,
            I => \N__47779\
        );

    \I__11445\ : SRMux
    port map (
            O => \N__48135\,
            I => \N__47779\
        );

    \I__11444\ : SRMux
    port map (
            O => \N__48134\,
            I => \N__47779\
        );

    \I__11443\ : SRMux
    port map (
            O => \N__48133\,
            I => \N__47779\
        );

    \I__11442\ : SRMux
    port map (
            O => \N__48132\,
            I => \N__47779\
        );

    \I__11441\ : SRMux
    port map (
            O => \N__48131\,
            I => \N__47779\
        );

    \I__11440\ : SRMux
    port map (
            O => \N__48130\,
            I => \N__47779\
        );

    \I__11439\ : SRMux
    port map (
            O => \N__48129\,
            I => \N__47779\
        );

    \I__11438\ : SRMux
    port map (
            O => \N__48128\,
            I => \N__47779\
        );

    \I__11437\ : SRMux
    port map (
            O => \N__48127\,
            I => \N__47779\
        );

    \I__11436\ : SRMux
    port map (
            O => \N__48126\,
            I => \N__47779\
        );

    \I__11435\ : SRMux
    port map (
            O => \N__48125\,
            I => \N__47779\
        );

    \I__11434\ : SRMux
    port map (
            O => \N__48124\,
            I => \N__47779\
        );

    \I__11433\ : SRMux
    port map (
            O => \N__48123\,
            I => \N__47779\
        );

    \I__11432\ : SRMux
    port map (
            O => \N__48122\,
            I => \N__47779\
        );

    \I__11431\ : SRMux
    port map (
            O => \N__48121\,
            I => \N__47779\
        );

    \I__11430\ : SRMux
    port map (
            O => \N__48120\,
            I => \N__47779\
        );

    \I__11429\ : SRMux
    port map (
            O => \N__48119\,
            I => \N__47779\
        );

    \I__11428\ : SRMux
    port map (
            O => \N__48118\,
            I => \N__47779\
        );

    \I__11427\ : SRMux
    port map (
            O => \N__48117\,
            I => \N__47779\
        );

    \I__11426\ : Glb2LocalMux
    port map (
            O => \N__48114\,
            I => \N__47779\
        );

    \I__11425\ : SRMux
    port map (
            O => \N__48113\,
            I => \N__47779\
        );

    \I__11424\ : SRMux
    port map (
            O => \N__48112\,
            I => \N__47779\
        );

    \I__11423\ : SRMux
    port map (
            O => \N__48111\,
            I => \N__47779\
        );

    \I__11422\ : SRMux
    port map (
            O => \N__48110\,
            I => \N__47779\
        );

    \I__11421\ : SRMux
    port map (
            O => \N__48109\,
            I => \N__47779\
        );

    \I__11420\ : SRMux
    port map (
            O => \N__48108\,
            I => \N__47779\
        );

    \I__11419\ : SRMux
    port map (
            O => \N__48107\,
            I => \N__47779\
        );

    \I__11418\ : SRMux
    port map (
            O => \N__48106\,
            I => \N__47779\
        );

    \I__11417\ : SRMux
    port map (
            O => \N__48105\,
            I => \N__47779\
        );

    \I__11416\ : SRMux
    port map (
            O => \N__48104\,
            I => \N__47779\
        );

    \I__11415\ : SRMux
    port map (
            O => \N__48103\,
            I => \N__47779\
        );

    \I__11414\ : SRMux
    port map (
            O => \N__48102\,
            I => \N__47779\
        );

    \I__11413\ : SRMux
    port map (
            O => \N__48101\,
            I => \N__47779\
        );

    \I__11412\ : SRMux
    port map (
            O => \N__48100\,
            I => \N__47779\
        );

    \I__11411\ : SRMux
    port map (
            O => \N__48099\,
            I => \N__47779\
        );

    \I__11410\ : SRMux
    port map (
            O => \N__48098\,
            I => \N__47779\
        );

    \I__11409\ : SRMux
    port map (
            O => \N__48097\,
            I => \N__47779\
        );

    \I__11408\ : SRMux
    port map (
            O => \N__48096\,
            I => \N__47779\
        );

    \I__11407\ : SRMux
    port map (
            O => \N__48095\,
            I => \N__47779\
        );

    \I__11406\ : SRMux
    port map (
            O => \N__48094\,
            I => \N__47779\
        );

    \I__11405\ : SRMux
    port map (
            O => \N__48093\,
            I => \N__47779\
        );

    \I__11404\ : SRMux
    port map (
            O => \N__48092\,
            I => \N__47779\
        );

    \I__11403\ : SRMux
    port map (
            O => \N__48091\,
            I => \N__47779\
        );

    \I__11402\ : SRMux
    port map (
            O => \N__48090\,
            I => \N__47779\
        );

    \I__11401\ : SRMux
    port map (
            O => \N__48089\,
            I => \N__47779\
        );

    \I__11400\ : SRMux
    port map (
            O => \N__48088\,
            I => \N__47779\
        );

    \I__11399\ : GlobalMux
    port map (
            O => \N__47779\,
            I => \N__47776\
        );

    \I__11398\ : gio2CtrlBuf
    port map (
            O => \N__47776\,
            I => red_c_g
        );

    \I__11397\ : CascadeMux
    port map (
            O => \N__47773\,
            I => \N__47768\
        );

    \I__11396\ : CascadeMux
    port map (
            O => \N__47772\,
            I => \N__47765\
        );

    \I__11395\ : InMux
    port map (
            O => \N__47771\,
            I => \N__47762\
        );

    \I__11394\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47757\
        );

    \I__11393\ : InMux
    port map (
            O => \N__47765\,
            I => \N__47757\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__47762\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__47757\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__11390\ : InMux
    port map (
            O => \N__47752\,
            I => \N__47749\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__47749\,
            I => \N__47746\
        );

    \I__11388\ : Span4Mux_v
    port map (
            O => \N__47746\,
            I => \N__47743\
        );

    \I__11387\ : Odrv4
    port map (
            O => \N__47743\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__11386\ : InMux
    port map (
            O => \N__47740\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__11385\ : CascadeMux
    port map (
            O => \N__47737\,
            I => \N__47732\
        );

    \I__11384\ : CascadeMux
    port map (
            O => \N__47736\,
            I => \N__47729\
        );

    \I__11383\ : InMux
    port map (
            O => \N__47735\,
            I => \N__47726\
        );

    \I__11382\ : InMux
    port map (
            O => \N__47732\,
            I => \N__47721\
        );

    \I__11381\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47721\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__47726\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__11379\ : LocalMux
    port map (
            O => \N__47721\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__11378\ : InMux
    port map (
            O => \N__47716\,
            I => \N__47713\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__47713\,
            I => \N__47710\
        );

    \I__11376\ : Span4Mux_v
    port map (
            O => \N__47710\,
            I => \N__47707\
        );

    \I__11375\ : Odrv4
    port map (
            O => \N__47707\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__11374\ : InMux
    port map (
            O => \N__47704\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__11373\ : InMux
    port map (
            O => \N__47701\,
            I => \N__47696\
        );

    \I__11372\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47691\
        );

    \I__11371\ : InMux
    port map (
            O => \N__47699\,
            I => \N__47691\
        );

    \I__11370\ : LocalMux
    port map (
            O => \N__47696\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__47691\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__11368\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47683\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__47683\,
            I => \N__47680\
        );

    \I__11366\ : Span4Mux_h
    port map (
            O => \N__47680\,
            I => \N__47677\
        );

    \I__11365\ : Odrv4
    port map (
            O => \N__47677\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__11364\ : InMux
    port map (
            O => \N__47674\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__11363\ : InMux
    port map (
            O => \N__47671\,
            I => \N__47666\
        );

    \I__11362\ : InMux
    port map (
            O => \N__47670\,
            I => \N__47661\
        );

    \I__11361\ : InMux
    port map (
            O => \N__47669\,
            I => \N__47661\
        );

    \I__11360\ : LocalMux
    port map (
            O => \N__47666\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__11359\ : LocalMux
    port map (
            O => \N__47661\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__11358\ : CascadeMux
    port map (
            O => \N__47656\,
            I => \N__47653\
        );

    \I__11357\ : InMux
    port map (
            O => \N__47653\,
            I => \N__47650\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__47650\,
            I => \N__47647\
        );

    \I__11355\ : Span4Mux_h
    port map (
            O => \N__47647\,
            I => \N__47644\
        );

    \I__11354\ : Odrv4
    port map (
            O => \N__47644\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__11353\ : InMux
    port map (
            O => \N__47641\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__11352\ : CascadeMux
    port map (
            O => \N__47638\,
            I => \N__47633\
        );

    \I__11351\ : CascadeMux
    port map (
            O => \N__47637\,
            I => \N__47630\
        );

    \I__11350\ : InMux
    port map (
            O => \N__47636\,
            I => \N__47627\
        );

    \I__11349\ : InMux
    port map (
            O => \N__47633\,
            I => \N__47622\
        );

    \I__11348\ : InMux
    port map (
            O => \N__47630\,
            I => \N__47622\
        );

    \I__11347\ : LocalMux
    port map (
            O => \N__47627\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__11346\ : LocalMux
    port map (
            O => \N__47622\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__11345\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47614\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__47614\,
            I => \N__47611\
        );

    \I__11343\ : Span4Mux_h
    port map (
            O => \N__47611\,
            I => \N__47608\
        );

    \I__11342\ : Odrv4
    port map (
            O => \N__47608\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__11341\ : InMux
    port map (
            O => \N__47605\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__11340\ : CascadeMux
    port map (
            O => \N__47602\,
            I => \N__47597\
        );

    \I__11339\ : CascadeMux
    port map (
            O => \N__47601\,
            I => \N__47594\
        );

    \I__11338\ : InMux
    port map (
            O => \N__47600\,
            I => \N__47591\
        );

    \I__11337\ : InMux
    port map (
            O => \N__47597\,
            I => \N__47586\
        );

    \I__11336\ : InMux
    port map (
            O => \N__47594\,
            I => \N__47586\
        );

    \I__11335\ : LocalMux
    port map (
            O => \N__47591\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__47586\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__11333\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47578\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__47578\,
            I => \N__47575\
        );

    \I__11331\ : Span4Mux_h
    port map (
            O => \N__47575\,
            I => \N__47572\
        );

    \I__11330\ : Odrv4
    port map (
            O => \N__47572\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__11329\ : InMux
    port map (
            O => \N__47569\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__11328\ : InMux
    port map (
            O => \N__47566\,
            I => \N__47561\
        );

    \I__11327\ : InMux
    port map (
            O => \N__47565\,
            I => \N__47558\
        );

    \I__11326\ : InMux
    port map (
            O => \N__47564\,
            I => \N__47555\
        );

    \I__11325\ : LocalMux
    port map (
            O => \N__47561\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__11324\ : LocalMux
    port map (
            O => \N__47558\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__47555\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__11322\ : InMux
    port map (
            O => \N__47548\,
            I => \N__47545\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__47545\,
            I => \N__47542\
        );

    \I__11320\ : Odrv4
    port map (
            O => \N__47542\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__11319\ : InMux
    port map (
            O => \N__47539\,
            I => \bfn_18_26_0_\
        );

    \I__11318\ : InMux
    port map (
            O => \N__47536\,
            I => \N__47531\
        );

    \I__11317\ : InMux
    port map (
            O => \N__47535\,
            I => \N__47528\
        );

    \I__11316\ : InMux
    port map (
            O => \N__47534\,
            I => \N__47525\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__47531\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__47528\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__47525\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__11312\ : CascadeMux
    port map (
            O => \N__47518\,
            I => \N__47515\
        );

    \I__11311\ : InMux
    port map (
            O => \N__47515\,
            I => \N__47512\
        );

    \I__11310\ : LocalMux
    port map (
            O => \N__47512\,
            I => \N__47509\
        );

    \I__11309\ : Odrv4
    port map (
            O => \N__47509\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__11308\ : InMux
    port map (
            O => \N__47506\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__11307\ : CascadeMux
    port map (
            O => \N__47503\,
            I => \N__47498\
        );

    \I__11306\ : CascadeMux
    port map (
            O => \N__47502\,
            I => \N__47495\
        );

    \I__11305\ : InMux
    port map (
            O => \N__47501\,
            I => \N__47492\
        );

    \I__11304\ : InMux
    port map (
            O => \N__47498\,
            I => \N__47487\
        );

    \I__11303\ : InMux
    port map (
            O => \N__47495\,
            I => \N__47487\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__47492\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__47487\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__11300\ : InMux
    port map (
            O => \N__47482\,
            I => \N__47478\
        );

    \I__11299\ : CascadeMux
    port map (
            O => \N__47481\,
            I => \N__47475\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__47478\,
            I => \N__47472\
        );

    \I__11297\ : InMux
    port map (
            O => \N__47475\,
            I => \N__47469\
        );

    \I__11296\ : Span4Mux_h
    port map (
            O => \N__47472\,
            I => \N__47466\
        );

    \I__11295\ : LocalMux
    port map (
            O => \N__47469\,
            I => \N__47463\
        );

    \I__11294\ : Span4Mux_v
    port map (
            O => \N__47466\,
            I => \N__47460\
        );

    \I__11293\ : Span4Mux_h
    port map (
            O => \N__47463\,
            I => \N__47457\
        );

    \I__11292\ : Odrv4
    port map (
            O => \N__47460\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__11291\ : Odrv4
    port map (
            O => \N__47457\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__11290\ : InMux
    port map (
            O => \N__47452\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__11289\ : CascadeMux
    port map (
            O => \N__47449\,
            I => \N__47444\
        );

    \I__11288\ : CascadeMux
    port map (
            O => \N__47448\,
            I => \N__47441\
        );

    \I__11287\ : InMux
    port map (
            O => \N__47447\,
            I => \N__47438\
        );

    \I__11286\ : InMux
    port map (
            O => \N__47444\,
            I => \N__47433\
        );

    \I__11285\ : InMux
    port map (
            O => \N__47441\,
            I => \N__47433\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__47438\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__11283\ : LocalMux
    port map (
            O => \N__47433\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__11282\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47422\
        );

    \I__11281\ : InMux
    port map (
            O => \N__47427\,
            I => \N__47419\
        );

    \I__11280\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47413\
        );

    \I__11279\ : InMux
    port map (
            O => \N__47425\,
            I => \N__47413\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__47422\,
            I => \N__47410\
        );

    \I__11277\ : LocalMux
    port map (
            O => \N__47419\,
            I => \N__47407\
        );

    \I__11276\ : InMux
    port map (
            O => \N__47418\,
            I => \N__47404\
        );

    \I__11275\ : LocalMux
    port map (
            O => \N__47413\,
            I => \N__47399\
        );

    \I__11274\ : Span4Mux_h
    port map (
            O => \N__47410\,
            I => \N__47399\
        );

    \I__11273\ : Span4Mux_h
    port map (
            O => \N__47407\,
            I => \N__47394\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47394\
        );

    \I__11271\ : Span4Mux_v
    port map (
            O => \N__47399\,
            I => \N__47391\
        );

    \I__11270\ : Span4Mux_h
    port map (
            O => \N__47394\,
            I => \N__47388\
        );

    \I__11269\ : Odrv4
    port map (
            O => \N__47391\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__11268\ : Odrv4
    port map (
            O => \N__47388\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__11267\ : InMux
    port map (
            O => \N__47383\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__11266\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47375\
        );

    \I__11265\ : InMux
    port map (
            O => \N__47379\,
            I => \N__47370\
        );

    \I__11264\ : InMux
    port map (
            O => \N__47378\,
            I => \N__47370\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__47375\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__11262\ : LocalMux
    port map (
            O => \N__47370\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__11261\ : InMux
    port map (
            O => \N__47365\,
            I => \N__47358\
        );

    \I__11260\ : CascadeMux
    port map (
            O => \N__47364\,
            I => \N__47355\
        );

    \I__11259\ : CascadeMux
    port map (
            O => \N__47363\,
            I => \N__47351\
        );

    \I__11258\ : InMux
    port map (
            O => \N__47362\,
            I => \N__47348\
        );

    \I__11257\ : InMux
    port map (
            O => \N__47361\,
            I => \N__47345\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__47358\,
            I => \N__47342\
        );

    \I__11255\ : InMux
    port map (
            O => \N__47355\,
            I => \N__47339\
        );

    \I__11254\ : InMux
    port map (
            O => \N__47354\,
            I => \N__47336\
        );

    \I__11253\ : InMux
    port map (
            O => \N__47351\,
            I => \N__47333\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__47348\,
            I => \N__47328\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__47345\,
            I => \N__47328\
        );

    \I__11250\ : Span4Mux_h
    port map (
            O => \N__47342\,
            I => \N__47319\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__47339\,
            I => \N__47319\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__47336\,
            I => \N__47319\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__47333\,
            I => \N__47319\
        );

    \I__11246\ : Span4Mux_v
    port map (
            O => \N__47328\,
            I => \N__47314\
        );

    \I__11245\ : Span4Mux_h
    port map (
            O => \N__47319\,
            I => \N__47314\
        );

    \I__11244\ : Odrv4
    port map (
            O => \N__47314\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__11243\ : InMux
    port map (
            O => \N__47311\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__11242\ : InMux
    port map (
            O => \N__47308\,
            I => \N__47303\
        );

    \I__11241\ : InMux
    port map (
            O => \N__47307\,
            I => \N__47298\
        );

    \I__11240\ : InMux
    port map (
            O => \N__47306\,
            I => \N__47298\
        );

    \I__11239\ : LocalMux
    port map (
            O => \N__47303\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__47298\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__11237\ : InMux
    port map (
            O => \N__47293\,
            I => \N__47290\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__47290\,
            I => \N__47286\
        );

    \I__11235\ : InMux
    port map (
            O => \N__47289\,
            I => \N__47283\
        );

    \I__11234\ : Span4Mux_v
    port map (
            O => \N__47286\,
            I => \N__47279\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__47283\,
            I => \N__47276\
        );

    \I__11232\ : InMux
    port map (
            O => \N__47282\,
            I => \N__47273\
        );

    \I__11231\ : Span4Mux_v
    port map (
            O => \N__47279\,
            I => \N__47268\
        );

    \I__11230\ : Span4Mux_v
    port map (
            O => \N__47276\,
            I => \N__47268\
        );

    \I__11229\ : LocalMux
    port map (
            O => \N__47273\,
            I => \N__47265\
        );

    \I__11228\ : Span4Mux_h
    port map (
            O => \N__47268\,
            I => \N__47262\
        );

    \I__11227\ : Odrv12
    port map (
            O => \N__47265\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__11226\ : Odrv4
    port map (
            O => \N__47262\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__11225\ : InMux
    port map (
            O => \N__47257\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__11224\ : CascadeMux
    port map (
            O => \N__47254\,
            I => \N__47249\
        );

    \I__11223\ : CascadeMux
    port map (
            O => \N__47253\,
            I => \N__47246\
        );

    \I__11222\ : InMux
    port map (
            O => \N__47252\,
            I => \N__47243\
        );

    \I__11221\ : InMux
    port map (
            O => \N__47249\,
            I => \N__47238\
        );

    \I__11220\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47238\
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__47243\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__11218\ : LocalMux
    port map (
            O => \N__47238\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__11217\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47229\
        );

    \I__11216\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47225\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47222\
        );

    \I__11214\ : InMux
    port map (
            O => \N__47228\,
            I => \N__47219\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__47225\,
            I => \N__47216\
        );

    \I__11212\ : Span12Mux_h
    port map (
            O => \N__47222\,
            I => \N__47211\
        );

    \I__11211\ : LocalMux
    port map (
            O => \N__47219\,
            I => \N__47211\
        );

    \I__11210\ : Span4Mux_h
    port map (
            O => \N__47216\,
            I => \N__47208\
        );

    \I__11209\ : Odrv12
    port map (
            O => \N__47211\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__11208\ : Odrv4
    port map (
            O => \N__47208\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__11207\ : InMux
    port map (
            O => \N__47203\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__11206\ : CascadeMux
    port map (
            O => \N__47200\,
            I => \N__47195\
        );

    \I__11205\ : CascadeMux
    port map (
            O => \N__47199\,
            I => \N__47192\
        );

    \I__11204\ : InMux
    port map (
            O => \N__47198\,
            I => \N__47189\
        );

    \I__11203\ : InMux
    port map (
            O => \N__47195\,
            I => \N__47184\
        );

    \I__11202\ : InMux
    port map (
            O => \N__47192\,
            I => \N__47184\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__47189\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__47184\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__11199\ : InMux
    port map (
            O => \N__47179\,
            I => \N__47176\
        );

    \I__11198\ : LocalMux
    port map (
            O => \N__47176\,
            I => \N__47173\
        );

    \I__11197\ : Span4Mux_h
    port map (
            O => \N__47173\,
            I => \N__47169\
        );

    \I__11196\ : InMux
    port map (
            O => \N__47172\,
            I => \N__47165\
        );

    \I__11195\ : Span4Mux_h
    port map (
            O => \N__47169\,
            I => \N__47162\
        );

    \I__11194\ : InMux
    port map (
            O => \N__47168\,
            I => \N__47159\
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__47165\,
            I => \N__47156\
        );

    \I__11192\ : Sp12to4
    port map (
            O => \N__47162\,
            I => \N__47151\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__47159\,
            I => \N__47151\
        );

    \I__11190\ : Span4Mux_h
    port map (
            O => \N__47156\,
            I => \N__47148\
        );

    \I__11189\ : Odrv12
    port map (
            O => \N__47151\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__11188\ : Odrv4
    port map (
            O => \N__47148\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__11187\ : InMux
    port map (
            O => \N__47143\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__11186\ : InMux
    port map (
            O => \N__47140\,
            I => \N__47135\
        );

    \I__11185\ : InMux
    port map (
            O => \N__47139\,
            I => \N__47132\
        );

    \I__11184\ : InMux
    port map (
            O => \N__47138\,
            I => \N__47129\
        );

    \I__11183\ : LocalMux
    port map (
            O => \N__47135\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__47132\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__47129\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__11180\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47119\
        );

    \I__11179\ : LocalMux
    port map (
            O => \N__47119\,
            I => \N__47114\
        );

    \I__11178\ : CascadeMux
    port map (
            O => \N__47118\,
            I => \N__47111\
        );

    \I__11177\ : CascadeMux
    port map (
            O => \N__47117\,
            I => \N__47108\
        );

    \I__11176\ : Span4Mux_h
    port map (
            O => \N__47114\,
            I => \N__47105\
        );

    \I__11175\ : InMux
    port map (
            O => \N__47111\,
            I => \N__47102\
        );

    \I__11174\ : InMux
    port map (
            O => \N__47108\,
            I => \N__47099\
        );

    \I__11173\ : Span4Mux_v
    port map (
            O => \N__47105\,
            I => \N__47096\
        );

    \I__11172\ : LocalMux
    port map (
            O => \N__47102\,
            I => \N__47093\
        );

    \I__11171\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47090\
        );

    \I__11170\ : Span4Mux_h
    port map (
            O => \N__47096\,
            I => \N__47087\
        );

    \I__11169\ : Span4Mux_v
    port map (
            O => \N__47093\,
            I => \N__47082\
        );

    \I__11168\ : Span4Mux_h
    port map (
            O => \N__47090\,
            I => \N__47082\
        );

    \I__11167\ : Odrv4
    port map (
            O => \N__47087\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__11166\ : Odrv4
    port map (
            O => \N__47082\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__11165\ : InMux
    port map (
            O => \N__47077\,
            I => \bfn_18_25_0_\
        );

    \I__11164\ : InMux
    port map (
            O => \N__47074\,
            I => \N__47069\
        );

    \I__11163\ : InMux
    port map (
            O => \N__47073\,
            I => \N__47066\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47072\,
            I => \N__47063\
        );

    \I__11161\ : LocalMux
    port map (
            O => \N__47069\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__11160\ : LocalMux
    port map (
            O => \N__47066\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__11159\ : LocalMux
    port map (
            O => \N__47063\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47056\,
            I => \N__47053\
        );

    \I__11157\ : LocalMux
    port map (
            O => \N__47053\,
            I => \N__47050\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__47050\,
            I => \N__47047\
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__47047\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__11154\ : InMux
    port map (
            O => \N__47044\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__11153\ : CascadeMux
    port map (
            O => \N__47041\,
            I => \N__47036\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__47040\,
            I => \N__47033\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47039\,
            I => \N__47030\
        );

    \I__11150\ : InMux
    port map (
            O => \N__47036\,
            I => \N__47025\
        );

    \I__11149\ : InMux
    port map (
            O => \N__47033\,
            I => \N__47025\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__47030\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__47025\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__11146\ : InMux
    port map (
            O => \N__47020\,
            I => \N__47015\
        );

    \I__11145\ : InMux
    port map (
            O => \N__47019\,
            I => \N__47012\
        );

    \I__11144\ : InMux
    port map (
            O => \N__47018\,
            I => \N__47009\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__47015\,
            I => \N__47002\
        );

    \I__11142\ : LocalMux
    port map (
            O => \N__47012\,
            I => \N__47002\
        );

    \I__11141\ : LocalMux
    port map (
            O => \N__47009\,
            I => \N__47002\
        );

    \I__11140\ : Span4Mux_h
    port map (
            O => \N__47002\,
            I => \N__46999\
        );

    \I__11139\ : Odrv4
    port map (
            O => \N__46999\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__11138\ : InMux
    port map (
            O => \N__46996\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__11137\ : InMux
    port map (
            O => \N__46993\,
            I => \N__46988\
        );

    \I__11136\ : InMux
    port map (
            O => \N__46992\,
            I => \N__46983\
        );

    \I__11135\ : InMux
    port map (
            O => \N__46991\,
            I => \N__46983\
        );

    \I__11134\ : LocalMux
    port map (
            O => \N__46988\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__11133\ : LocalMux
    port map (
            O => \N__46983\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__11132\ : InMux
    port map (
            O => \N__46978\,
            I => \N__46975\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__46975\,
            I => \N__46972\
        );

    \I__11130\ : Span4Mux_v
    port map (
            O => \N__46972\,
            I => \N__46967\
        );

    \I__11129\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46964\
        );

    \I__11128\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46961\
        );

    \I__11127\ : Span4Mux_v
    port map (
            O => \N__46967\,
            I => \N__46958\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__46964\,
            I => \N__46953\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__46961\,
            I => \N__46953\
        );

    \I__11124\ : Span4Mux_h
    port map (
            O => \N__46958\,
            I => \N__46950\
        );

    \I__11123\ : Span4Mux_h
    port map (
            O => \N__46953\,
            I => \N__46947\
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__46950\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__11121\ : Odrv4
    port map (
            O => \N__46947\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__11120\ : InMux
    port map (
            O => \N__46942\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__11119\ : InMux
    port map (
            O => \N__46939\,
            I => \N__46934\
        );

    \I__11118\ : InMux
    port map (
            O => \N__46938\,
            I => \N__46929\
        );

    \I__11117\ : InMux
    port map (
            O => \N__46937\,
            I => \N__46929\
        );

    \I__11116\ : LocalMux
    port map (
            O => \N__46934\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__46929\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__11114\ : InMux
    port map (
            O => \N__46924\,
            I => \N__46921\
        );

    \I__11113\ : LocalMux
    port map (
            O => \N__46921\,
            I => \N__46918\
        );

    \I__11112\ : Span4Mux_h
    port map (
            O => \N__46918\,
            I => \N__46913\
        );

    \I__11111\ : InMux
    port map (
            O => \N__46917\,
            I => \N__46910\
        );

    \I__11110\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46907\
        );

    \I__11109\ : Span4Mux_h
    port map (
            O => \N__46913\,
            I => \N__46904\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__46910\,
            I => \N__46899\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__46907\,
            I => \N__46899\
        );

    \I__11106\ : Span4Mux_v
    port map (
            O => \N__46904\,
            I => \N__46896\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__46899\,
            I => \N__46893\
        );

    \I__11104\ : Odrv4
    port map (
            O => \N__46896\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__11103\ : Odrv4
    port map (
            O => \N__46893\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__11102\ : InMux
    port map (
            O => \N__46888\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__11101\ : CascadeMux
    port map (
            O => \N__46885\,
            I => \N__46880\
        );

    \I__11100\ : CascadeMux
    port map (
            O => \N__46884\,
            I => \N__46877\
        );

    \I__11099\ : InMux
    port map (
            O => \N__46883\,
            I => \N__46874\
        );

    \I__11098\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46869\
        );

    \I__11097\ : InMux
    port map (
            O => \N__46877\,
            I => \N__46869\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__46874\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__11095\ : LocalMux
    port map (
            O => \N__46869\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__11094\ : CascadeMux
    port map (
            O => \N__46864\,
            I => \N__46861\
        );

    \I__11093\ : InMux
    port map (
            O => \N__46861\,
            I => \N__46857\
        );

    \I__11092\ : CascadeMux
    port map (
            O => \N__46860\,
            I => \N__46853\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__46857\,
            I => \N__46849\
        );

    \I__11090\ : InMux
    port map (
            O => \N__46856\,
            I => \N__46846\
        );

    \I__11089\ : InMux
    port map (
            O => \N__46853\,
            I => \N__46843\
        );

    \I__11088\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46840\
        );

    \I__11087\ : Span4Mux_h
    port map (
            O => \N__46849\,
            I => \N__46837\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__46846\,
            I => \N__46834\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__46843\,
            I => \N__46831\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__46840\,
            I => \N__46828\
        );

    \I__11083\ : Span4Mux_v
    port map (
            O => \N__46837\,
            I => \N__46825\
        );

    \I__11082\ : Span4Mux_v
    port map (
            O => \N__46834\,
            I => \N__46818\
        );

    \I__11081\ : Span4Mux_v
    port map (
            O => \N__46831\,
            I => \N__46818\
        );

    \I__11080\ : Span4Mux_h
    port map (
            O => \N__46828\,
            I => \N__46818\
        );

    \I__11079\ : Odrv4
    port map (
            O => \N__46825\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__46818\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__11077\ : InMux
    port map (
            O => \N__46813\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__11076\ : CascadeMux
    port map (
            O => \N__46810\,
            I => \N__46805\
        );

    \I__11075\ : CascadeMux
    port map (
            O => \N__46809\,
            I => \N__46802\
        );

    \I__11074\ : InMux
    port map (
            O => \N__46808\,
            I => \N__46799\
        );

    \I__11073\ : InMux
    port map (
            O => \N__46805\,
            I => \N__46794\
        );

    \I__11072\ : InMux
    port map (
            O => \N__46802\,
            I => \N__46794\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__46799\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__46794\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__11069\ : InMux
    port map (
            O => \N__46789\,
            I => \N__46785\
        );

    \I__11068\ : InMux
    port map (
            O => \N__46788\,
            I => \N__46782\
        );

    \I__11067\ : LocalMux
    port map (
            O => \N__46785\,
            I => \N__46779\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__46782\,
            I => \N__46776\
        );

    \I__11065\ : Span12Mux_v
    port map (
            O => \N__46779\,
            I => \N__46773\
        );

    \I__11064\ : Span4Mux_h
    port map (
            O => \N__46776\,
            I => \N__46770\
        );

    \I__11063\ : Odrv12
    port map (
            O => \N__46773\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__11062\ : Odrv4
    port map (
            O => \N__46770\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__11061\ : InMux
    port map (
            O => \N__46765\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__11060\ : InMux
    port map (
            O => \N__46762\,
            I => \N__46757\
        );

    \I__11059\ : InMux
    port map (
            O => \N__46761\,
            I => \N__46754\
        );

    \I__11058\ : InMux
    port map (
            O => \N__46760\,
            I => \N__46751\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__46757\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__46754\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__46751\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__11054\ : InMux
    port map (
            O => \N__46744\,
            I => \N__46741\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__46741\,
            I => \N__46737\
        );

    \I__11052\ : InMux
    port map (
            O => \N__46740\,
            I => \N__46734\
        );

    \I__11051\ : Span4Mux_v
    port map (
            O => \N__46737\,
            I => \N__46731\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__46734\,
            I => \N__46728\
        );

    \I__11049\ : Span4Mux_h
    port map (
            O => \N__46731\,
            I => \N__46725\
        );

    \I__11048\ : Span4Mux_h
    port map (
            O => \N__46728\,
            I => \N__46722\
        );

    \I__11047\ : Odrv4
    port map (
            O => \N__46725\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__11046\ : Odrv4
    port map (
            O => \N__46722\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__11045\ : InMux
    port map (
            O => \N__46717\,
            I => \bfn_18_24_0_\
        );

    \I__11044\ : InMux
    port map (
            O => \N__46714\,
            I => \N__46709\
        );

    \I__11043\ : InMux
    port map (
            O => \N__46713\,
            I => \N__46706\
        );

    \I__11042\ : InMux
    port map (
            O => \N__46712\,
            I => \N__46703\
        );

    \I__11041\ : LocalMux
    port map (
            O => \N__46709\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__46706\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__46703\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__11038\ : InMux
    port map (
            O => \N__46696\,
            I => \N__46693\
        );

    \I__11037\ : LocalMux
    port map (
            O => \N__46693\,
            I => \N__46689\
        );

    \I__11036\ : InMux
    port map (
            O => \N__46692\,
            I => \N__46686\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__46689\,
            I => \N__46683\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__46686\,
            I => \N__46680\
        );

    \I__11033\ : Span4Mux_h
    port map (
            O => \N__46683\,
            I => \N__46677\
        );

    \I__11032\ : Span4Mux_h
    port map (
            O => \N__46680\,
            I => \N__46674\
        );

    \I__11031\ : Odrv4
    port map (
            O => \N__46677\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__11030\ : Odrv4
    port map (
            O => \N__46674\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__11029\ : InMux
    port map (
            O => \N__46669\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__11028\ : CascadeMux
    port map (
            O => \N__46666\,
            I => \N__46663\
        );

    \I__11027\ : InMux
    port map (
            O => \N__46663\,
            I => \N__46660\
        );

    \I__11026\ : LocalMux
    port map (
            O => \N__46660\,
            I => \N__46657\
        );

    \I__11025\ : Span4Mux_h
    port map (
            O => \N__46657\,
            I => \N__46654\
        );

    \I__11024\ : Span4Mux_v
    port map (
            O => \N__46654\,
            I => \N__46651\
        );

    \I__11023\ : Odrv4
    port map (
            O => \N__46651\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__11022\ : CEMux
    port map (
            O => \N__46648\,
            I => \N__46645\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__46645\,
            I => \N__46638\
        );

    \I__11020\ : CEMux
    port map (
            O => \N__46644\,
            I => \N__46635\
        );

    \I__11019\ : CEMux
    port map (
            O => \N__46643\,
            I => \N__46632\
        );

    \I__11018\ : CEMux
    port map (
            O => \N__46642\,
            I => \N__46629\
        );

    \I__11017\ : CEMux
    port map (
            O => \N__46641\,
            I => \N__46625\
        );

    \I__11016\ : Span4Mux_v
    port map (
            O => \N__46638\,
            I => \N__46622\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__46635\,
            I => \N__46619\
        );

    \I__11014\ : LocalMux
    port map (
            O => \N__46632\,
            I => \N__46616\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__46629\,
            I => \N__46613\
        );

    \I__11012\ : CEMux
    port map (
            O => \N__46628\,
            I => \N__46610\
        );

    \I__11011\ : LocalMux
    port map (
            O => \N__46625\,
            I => \N__46607\
        );

    \I__11010\ : Span4Mux_v
    port map (
            O => \N__46622\,
            I => \N__46604\
        );

    \I__11009\ : Span4Mux_v
    port map (
            O => \N__46619\,
            I => \N__46601\
        );

    \I__11008\ : Span4Mux_v
    port map (
            O => \N__46616\,
            I => \N__46598\
        );

    \I__11007\ : Span4Mux_v
    port map (
            O => \N__46613\,
            I => \N__46593\
        );

    \I__11006\ : LocalMux
    port map (
            O => \N__46610\,
            I => \N__46593\
        );

    \I__11005\ : Span4Mux_h
    port map (
            O => \N__46607\,
            I => \N__46590\
        );

    \I__11004\ : Sp12to4
    port map (
            O => \N__46604\,
            I => \N__46583\
        );

    \I__11003\ : Sp12to4
    port map (
            O => \N__46601\,
            I => \N__46583\
        );

    \I__11002\ : Sp12to4
    port map (
            O => \N__46598\,
            I => \N__46583\
        );

    \I__11001\ : Span4Mux_v
    port map (
            O => \N__46593\,
            I => \N__46580\
        );

    \I__11000\ : Span4Mux_h
    port map (
            O => \N__46590\,
            I => \N__46577\
        );

    \I__10999\ : Odrv12
    port map (
            O => \N__46583\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10998\ : Odrv4
    port map (
            O => \N__46580\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10997\ : Odrv4
    port map (
            O => \N__46577\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10996\ : CascadeMux
    port map (
            O => \N__46570\,
            I => \N__46566\
        );

    \I__10995\ : InMux
    port map (
            O => \N__46569\,
            I => \N__46563\
        );

    \I__10994\ : InMux
    port map (
            O => \N__46566\,
            I => \N__46560\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__46563\,
            I => \N__46556\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__46560\,
            I => \N__46553\
        );

    \I__10991\ : CascadeMux
    port map (
            O => \N__46559\,
            I => \N__46550\
        );

    \I__10990\ : Span4Mux_h
    port map (
            O => \N__46556\,
            I => \N__46547\
        );

    \I__10989\ : Span12Mux_v
    port map (
            O => \N__46553\,
            I => \N__46544\
        );

    \I__10988\ : InMux
    port map (
            O => \N__46550\,
            I => \N__46541\
        );

    \I__10987\ : Span4Mux_h
    port map (
            O => \N__46547\,
            I => \N__46538\
        );

    \I__10986\ : Odrv12
    port map (
            O => \N__46544\,
            I => measured_delay_tr_4
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__46541\,
            I => measured_delay_tr_4
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__46538\,
            I => measured_delay_tr_4
        );

    \I__10983\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46528\
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__46528\,
            I => \N__46523\
        );

    \I__10981\ : InMux
    port map (
            O => \N__46527\,
            I => \N__46520\
        );

    \I__10980\ : InMux
    port map (
            O => \N__46526\,
            I => \N__46517\
        );

    \I__10979\ : Span4Mux_h
    port map (
            O => \N__46523\,
            I => \N__46513\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__46520\,
            I => \N__46510\
        );

    \I__10977\ : LocalMux
    port map (
            O => \N__46517\,
            I => \N__46507\
        );

    \I__10976\ : InMux
    port map (
            O => \N__46516\,
            I => \N__46504\
        );

    \I__10975\ : Span4Mux_h
    port map (
            O => \N__46513\,
            I => \N__46498\
        );

    \I__10974\ : Span4Mux_h
    port map (
            O => \N__46510\,
            I => \N__46491\
        );

    \I__10973\ : Span4Mux_v
    port map (
            O => \N__46507\,
            I => \N__46491\
        );

    \I__10972\ : LocalMux
    port map (
            O => \N__46504\,
            I => \N__46491\
        );

    \I__10971\ : InMux
    port map (
            O => \N__46503\,
            I => \N__46486\
        );

    \I__10970\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46486\
        );

    \I__10969\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46483\
        );

    \I__10968\ : Odrv4
    port map (
            O => \N__46498\,
            I => \delay_measurement_inst.N_425\
        );

    \I__10967\ : Odrv4
    port map (
            O => \N__46491\,
            I => \delay_measurement_inst.N_425\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__46486\,
            I => \delay_measurement_inst.N_425\
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__46483\,
            I => \delay_measurement_inst.N_425\
        );

    \I__10964\ : InMux
    port map (
            O => \N__46474\,
            I => \N__46470\
        );

    \I__10963\ : InMux
    port map (
            O => \N__46473\,
            I => \N__46467\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__46470\,
            I => \N__46464\
        );

    \I__10961\ : LocalMux
    port map (
            O => \N__46467\,
            I => \N__46460\
        );

    \I__10960\ : Span4Mux_h
    port map (
            O => \N__46464\,
            I => \N__46457\
        );

    \I__10959\ : InMux
    port map (
            O => \N__46463\,
            I => \N__46454\
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__46460\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10957\ : Odrv4
    port map (
            O => \N__46457\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10956\ : LocalMux
    port map (
            O => \N__46454\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__10955\ : InMux
    port map (
            O => \N__46447\,
            I => \N__46443\
        );

    \I__10954\ : InMux
    port map (
            O => \N__46446\,
            I => \N__46440\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__46443\,
            I => \N__46433\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__46440\,
            I => \N__46433\
        );

    \I__10951\ : InMux
    port map (
            O => \N__46439\,
            I => \N__46430\
        );

    \I__10950\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46427\
        );

    \I__10949\ : Span4Mux_v
    port map (
            O => \N__46433\,
            I => \N__46424\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__46430\,
            I => \N__46419\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__46427\,
            I => \N__46419\
        );

    \I__10946\ : Span4Mux_h
    port map (
            O => \N__46424\,
            I => \N__46412\
        );

    \I__10945\ : Span4Mux_v
    port map (
            O => \N__46419\,
            I => \N__46409\
        );

    \I__10944\ : InMux
    port map (
            O => \N__46418\,
            I => \N__46402\
        );

    \I__10943\ : InMux
    port map (
            O => \N__46417\,
            I => \N__46402\
        );

    \I__10942\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46402\
        );

    \I__10941\ : InMux
    port map (
            O => \N__46415\,
            I => \N__46399\
        );

    \I__10940\ : Odrv4
    port map (
            O => \N__46412\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__10939\ : Odrv4
    port map (
            O => \N__46409\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__10938\ : LocalMux
    port map (
            O => \N__46402\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__46399\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__10936\ : InMux
    port map (
            O => \N__46390\,
            I => \N__46387\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__46387\,
            I => \N__46383\
        );

    \I__10934\ : InMux
    port map (
            O => \N__46386\,
            I => \N__46379\
        );

    \I__10933\ : Span4Mux_h
    port map (
            O => \N__46383\,
            I => \N__46376\
        );

    \I__10932\ : InMux
    port map (
            O => \N__46382\,
            I => \N__46373\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__46379\,
            I => \N__46370\
        );

    \I__10930\ : Span4Mux_v
    port map (
            O => \N__46376\,
            I => \N__46367\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__46373\,
            I => \N__46364\
        );

    \I__10928\ : Span4Mux_h
    port map (
            O => \N__46370\,
            I => \N__46361\
        );

    \I__10927\ : Odrv4
    port map (
            O => \N__46367\,
            I => measured_delay_tr_2
        );

    \I__10926\ : Odrv12
    port map (
            O => \N__46364\,
            I => measured_delay_tr_2
        );

    \I__10925\ : Odrv4
    port map (
            O => \N__46361\,
            I => measured_delay_tr_2
        );

    \I__10924\ : CEMux
    port map (
            O => \N__46354\,
            I => \N__46351\
        );

    \I__10923\ : LocalMux
    port map (
            O => \N__46351\,
            I => \N__46346\
        );

    \I__10922\ : CEMux
    port map (
            O => \N__46350\,
            I => \N__46340\
        );

    \I__10921\ : CEMux
    port map (
            O => \N__46349\,
            I => \N__46337\
        );

    \I__10920\ : Span4Mux_v
    port map (
            O => \N__46346\,
            I => \N__46334\
        );

    \I__10919\ : CEMux
    port map (
            O => \N__46345\,
            I => \N__46331\
        );

    \I__10918\ : CEMux
    port map (
            O => \N__46344\,
            I => \N__46328\
        );

    \I__10917\ : CEMux
    port map (
            O => \N__46343\,
            I => \N__46325\
        );

    \I__10916\ : LocalMux
    port map (
            O => \N__46340\,
            I => \N__46322\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__46337\,
            I => \N__46319\
        );

    \I__10914\ : Span4Mux_h
    port map (
            O => \N__46334\,
            I => \N__46314\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__46331\,
            I => \N__46314\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__46328\,
            I => \N__46311\
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__46325\,
            I => \N__46308\
        );

    \I__10910\ : Span4Mux_v
    port map (
            O => \N__46322\,
            I => \N__46305\
        );

    \I__10909\ : Span4Mux_v
    port map (
            O => \N__46319\,
            I => \N__46302\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__46314\,
            I => \N__46297\
        );

    \I__10907\ : Span4Mux_h
    port map (
            O => \N__46311\,
            I => \N__46297\
        );

    \I__10906\ : Span4Mux_h
    port map (
            O => \N__46308\,
            I => \N__46294\
        );

    \I__10905\ : Odrv4
    port map (
            O => \N__46305\,
            I => \delay_measurement_inst.N_280_i_0\
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__46302\,
            I => \delay_measurement_inst.N_280_i_0\
        );

    \I__10903\ : Odrv4
    port map (
            O => \N__46297\,
            I => \delay_measurement_inst.N_280_i_0\
        );

    \I__10902\ : Odrv4
    port map (
            O => \N__46294\,
            I => \delay_measurement_inst.N_280_i_0\
        );

    \I__10901\ : InMux
    port map (
            O => \N__46285\,
            I => \N__46279\
        );

    \I__10900\ : InMux
    port map (
            O => \N__46284\,
            I => \N__46279\
        );

    \I__10899\ : LocalMux
    port map (
            O => \N__46279\,
            I => \N__46276\
        );

    \I__10898\ : Span4Mux_h
    port map (
            O => \N__46276\,
            I => \N__46273\
        );

    \I__10897\ : Odrv4
    port map (
            O => \N__46273\,
            I => \delay_measurement_inst.N_286_1\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46265\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46262\
        );

    \I__10894\ : InMux
    port map (
            O => \N__46268\,
            I => \N__46259\
        );

    \I__10893\ : LocalMux
    port map (
            O => \N__46265\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__46262\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__46259\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__10890\ : InMux
    port map (
            O => \N__46252\,
            I => \N__46245\
        );

    \I__10889\ : InMux
    port map (
            O => \N__46251\,
            I => \N__46245\
        );

    \I__10888\ : InMux
    port map (
            O => \N__46250\,
            I => \N__46242\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46245\,
            I => \N__46235\
        );

    \I__10886\ : LocalMux
    port map (
            O => \N__46242\,
            I => \N__46232\
        );

    \I__10885\ : InMux
    port map (
            O => \N__46241\,
            I => \N__46229\
        );

    \I__10884\ : InMux
    port map (
            O => \N__46240\,
            I => \N__46226\
        );

    \I__10883\ : InMux
    port map (
            O => \N__46239\,
            I => \N__46221\
        );

    \I__10882\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46221\
        );

    \I__10881\ : Span4Mux_h
    port map (
            O => \N__46235\,
            I => \N__46216\
        );

    \I__10880\ : Span4Mux_v
    port map (
            O => \N__46232\,
            I => \N__46213\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__46229\,
            I => \N__46210\
        );

    \I__10878\ : LocalMux
    port map (
            O => \N__46226\,
            I => \N__46205\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46221\,
            I => \N__46205\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46220\,
            I => \N__46202\
        );

    \I__10875\ : InMux
    port map (
            O => \N__46219\,
            I => \N__46199\
        );

    \I__10874\ : Span4Mux_v
    port map (
            O => \N__46216\,
            I => \N__46196\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__46213\,
            I => \N__46191\
        );

    \I__10872\ : Span4Mux_v
    port map (
            O => \N__46210\,
            I => \N__46191\
        );

    \I__10871\ : Span12Mux_h
    port map (
            O => \N__46205\,
            I => \N__46184\
        );

    \I__10870\ : LocalMux
    port map (
            O => \N__46202\,
            I => \N__46184\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__46199\,
            I => \N__46184\
        );

    \I__10868\ : Odrv4
    port map (
            O => \N__46196\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__10867\ : Odrv4
    port map (
            O => \N__46191\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__10866\ : Odrv12
    port map (
            O => \N__46184\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__10865\ : CascadeMux
    port map (
            O => \N__46177\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16_cascade_\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46174\,
            I => \N__46171\
        );

    \I__10863\ : LocalMux
    port map (
            O => \N__46171\,
            I => \delay_measurement_inst.delay_tr_timer.N_415\
        );

    \I__10862\ : CascadeMux
    port map (
            O => \N__46168\,
            I => \N__46162\
        );

    \I__10861\ : CascadeMux
    port map (
            O => \N__46167\,
            I => \N__46159\
        );

    \I__10860\ : CascadeMux
    port map (
            O => \N__46166\,
            I => \N__46156\
        );

    \I__10859\ : InMux
    port map (
            O => \N__46165\,
            I => \N__46148\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46162\,
            I => \N__46148\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46145\
        );

    \I__10856\ : InMux
    port map (
            O => \N__46156\,
            I => \N__46142\
        );

    \I__10855\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46139\
        );

    \I__10854\ : InMux
    port map (
            O => \N__46154\,
            I => \N__46136\
        );

    \I__10853\ : CascadeMux
    port map (
            O => \N__46153\,
            I => \N__46132\
        );

    \I__10852\ : LocalMux
    port map (
            O => \N__46148\,
            I => \N__46129\
        );

    \I__10851\ : LocalMux
    port map (
            O => \N__46145\,
            I => \N__46122\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__46142\,
            I => \N__46122\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46139\,
            I => \N__46122\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46136\,
            I => \N__46119\
        );

    \I__10847\ : CascadeMux
    port map (
            O => \N__46135\,
            I => \N__46116\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46113\
        );

    \I__10845\ : Span4Mux_v
    port map (
            O => \N__46129\,
            I => \N__46108\
        );

    \I__10844\ : Span4Mux_v
    port map (
            O => \N__46122\,
            I => \N__46108\
        );

    \I__10843\ : Span4Mux_h
    port map (
            O => \N__46119\,
            I => \N__46105\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46116\,
            I => \N__46102\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46113\,
            I => \N__46099\
        );

    \I__10840\ : Span4Mux_h
    port map (
            O => \N__46108\,
            I => \N__46094\
        );

    \I__10839\ : Span4Mux_v
    port map (
            O => \N__46105\,
            I => \N__46094\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46102\,
            I => \delay_measurement_inst.N_373\
        );

    \I__10837\ : Odrv4
    port map (
            O => \N__46099\,
            I => \delay_measurement_inst.N_373\
        );

    \I__10836\ : Odrv4
    port map (
            O => \N__46094\,
            I => \delay_measurement_inst.N_373\
        );

    \I__10835\ : InMux
    port map (
            O => \N__46087\,
            I => \N__46083\
        );

    \I__10834\ : CascadeMux
    port map (
            O => \N__46086\,
            I => \N__46080\
        );

    \I__10833\ : LocalMux
    port map (
            O => \N__46083\,
            I => \N__46076\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46080\,
            I => \N__46073\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46079\,
            I => \N__46070\
        );

    \I__10830\ : Span4Mux_h
    port map (
            O => \N__46076\,
            I => \N__46065\
        );

    \I__10829\ : LocalMux
    port map (
            O => \N__46073\,
            I => \N__46065\
        );

    \I__10828\ : LocalMux
    port map (
            O => \N__46070\,
            I => \N__46062\
        );

    \I__10827\ : Span4Mux_h
    port map (
            O => \N__46065\,
            I => \N__46059\
        );

    \I__10826\ : Span4Mux_h
    port map (
            O => \N__46062\,
            I => \N__46056\
        );

    \I__10825\ : Odrv4
    port map (
            O => \N__46059\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__10824\ : Odrv4
    port map (
            O => \N__46056\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46051\,
            I => \N__46048\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46048\,
            I => \N__46043\
        );

    \I__10821\ : InMux
    port map (
            O => \N__46047\,
            I => \N__46040\
        );

    \I__10820\ : InMux
    port map (
            O => \N__46046\,
            I => \N__46037\
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__46043\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__46040\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10817\ : LocalMux
    port map (
            O => \N__46037\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46030\,
            I => \N__46025\
        );

    \I__10815\ : InMux
    port map (
            O => \N__46029\,
            I => \N__46022\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46028\,
            I => \N__46019\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46025\,
            I => \N__46016\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__46022\,
            I => \N__46013\
        );

    \I__10811\ : LocalMux
    port map (
            O => \N__46019\,
            I => \N__46010\
        );

    \I__10810\ : Span4Mux_h
    port map (
            O => \N__46016\,
            I => \N__46007\
        );

    \I__10809\ : Span4Mux_h
    port map (
            O => \N__46013\,
            I => \N__46004\
        );

    \I__10808\ : Odrv12
    port map (
            O => \N__46010\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10807\ : Odrv4
    port map (
            O => \N__46007\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10806\ : Odrv4
    port map (
            O => \N__46004\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__10805\ : InMux
    port map (
            O => \N__45997\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__10804\ : CascadeMux
    port map (
            O => \N__45994\,
            I => \N__45989\
        );

    \I__10803\ : CascadeMux
    port map (
            O => \N__45993\,
            I => \N__45986\
        );

    \I__10802\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45983\
        );

    \I__10801\ : InMux
    port map (
            O => \N__45989\,
            I => \N__45978\
        );

    \I__10800\ : InMux
    port map (
            O => \N__45986\,
            I => \N__45978\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__45983\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__45978\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__10797\ : CascadeMux
    port map (
            O => \N__45973\,
            I => \N__45970\
        );

    \I__10796\ : InMux
    port map (
            O => \N__45970\,
            I => \N__45965\
        );

    \I__10795\ : InMux
    port map (
            O => \N__45969\,
            I => \N__45962\
        );

    \I__10794\ : InMux
    port map (
            O => \N__45968\,
            I => \N__45959\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45954\
        );

    \I__10792\ : LocalMux
    port map (
            O => \N__45962\,
            I => \N__45954\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__45959\,
            I => \N__45951\
        );

    \I__10790\ : Span4Mux_h
    port map (
            O => \N__45954\,
            I => \N__45948\
        );

    \I__10789\ : Span4Mux_h
    port map (
            O => \N__45951\,
            I => \N__45945\
        );

    \I__10788\ : Odrv4
    port map (
            O => \N__45948\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__10787\ : Odrv4
    port map (
            O => \N__45945\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__10786\ : InMux
    port map (
            O => \N__45940\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__10785\ : InMux
    port map (
            O => \N__45937\,
            I => \N__45934\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__45934\,
            I => \N__45931\
        );

    \I__10783\ : Span4Mux_v
    port map (
            O => \N__45931\,
            I => \N__45927\
        );

    \I__10782\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45924\
        );

    \I__10781\ : Sp12to4
    port map (
            O => \N__45927\,
            I => \N__45917\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__45924\,
            I => \N__45917\
        );

    \I__10779\ : InMux
    port map (
            O => \N__45923\,
            I => \N__45914\
        );

    \I__10778\ : InMux
    port map (
            O => \N__45922\,
            I => \N__45911\
        );

    \I__10777\ : Odrv12
    port map (
            O => \N__45917\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__10776\ : LocalMux
    port map (
            O => \N__45914\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__45911\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__10774\ : InMux
    port map (
            O => \N__45904\,
            I => \N__45901\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__45901\,
            I => \N__45897\
        );

    \I__10772\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45893\
        );

    \I__10771\ : Span4Mux_h
    port map (
            O => \N__45897\,
            I => \N__45890\
        );

    \I__10770\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45887\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__45893\,
            I => \N__45884\
        );

    \I__10768\ : Odrv4
    port map (
            O => \N__45890\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__45887\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__10766\ : Odrv4
    port map (
            O => \N__45884\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__10765\ : CascadeMux
    port map (
            O => \N__45877\,
            I => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_\
        );

    \I__10764\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45867\
        );

    \I__10763\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45862\
        );

    \I__10762\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45862\
        );

    \I__10761\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45858\
        );

    \I__10760\ : InMux
    port map (
            O => \N__45870\,
            I => \N__45855\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__45867\,
            I => \N__45852\
        );

    \I__10758\ : LocalMux
    port map (
            O => \N__45862\,
            I => \N__45849\
        );

    \I__10757\ : InMux
    port map (
            O => \N__45861\,
            I => \N__45846\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__45858\,
            I => \N__45841\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__45855\,
            I => \N__45841\
        );

    \I__10754\ : Span4Mux_h
    port map (
            O => \N__45852\,
            I => \N__45838\
        );

    \I__10753\ : Span4Mux_v
    port map (
            O => \N__45849\,
            I => \N__45833\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__45846\,
            I => \N__45833\
        );

    \I__10751\ : Span4Mux_h
    port map (
            O => \N__45841\,
            I => \N__45830\
        );

    \I__10750\ : Odrv4
    port map (
            O => \N__45838\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10749\ : Odrv4
    port map (
            O => \N__45833\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10748\ : Odrv4
    port map (
            O => \N__45830\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__10747\ : CascadeMux
    port map (
            O => \N__45823\,
            I => \N__45819\
        );

    \I__10746\ : InMux
    port map (
            O => \N__45822\,
            I => \N__45815\
        );

    \I__10745\ : InMux
    port map (
            O => \N__45819\,
            I => \N__45812\
        );

    \I__10744\ : InMux
    port map (
            O => \N__45818\,
            I => \N__45809\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__45815\,
            I => \N__45802\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__45812\,
            I => \N__45802\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__45809\,
            I => \N__45802\
        );

    \I__10740\ : Span4Mux_v
    port map (
            O => \N__45802\,
            I => \N__45799\
        );

    \I__10739\ : Odrv4
    port map (
            O => \N__45799\,
            I => \il_max_comp2_D2\
        );

    \I__10738\ : InMux
    port map (
            O => \N__45796\,
            I => \N__45793\
        );

    \I__10737\ : LocalMux
    port map (
            O => \N__45793\,
            I => \N__45790\
        );

    \I__10736\ : Odrv12
    port map (
            O => \N__45790\,
            I => \phase_controller_slave.N_213\
        );

    \I__10735\ : InMux
    port map (
            O => \N__45787\,
            I => \N__45784\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__45784\,
            I => \N__45781\
        );

    \I__10733\ : Odrv12
    port map (
            O => \N__45781\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__10732\ : InMux
    port map (
            O => \N__45778\,
            I => \N__45775\
        );

    \I__10731\ : LocalMux
    port map (
            O => \N__45775\,
            I => \N__45771\
        );

    \I__10730\ : InMux
    port map (
            O => \N__45774\,
            I => \N__45768\
        );

    \I__10729\ : Span4Mux_h
    port map (
            O => \N__45771\,
            I => \N__45763\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__45768\,
            I => \N__45763\
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__45763\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__10726\ : InMux
    port map (
            O => \N__45760\,
            I => \N__45753\
        );

    \I__10725\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45750\
        );

    \I__10724\ : InMux
    port map (
            O => \N__45758\,
            I => \N__45747\
        );

    \I__10723\ : InMux
    port map (
            O => \N__45757\,
            I => \N__45744\
        );

    \I__10722\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45741\
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__45753\,
            I => \N__45736\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45736\
        );

    \I__10719\ : LocalMux
    port map (
            O => \N__45747\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45744\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__45741\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__10716\ : Odrv4
    port map (
            O => \N__45736\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__10715\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45723\
        );

    \I__10714\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45720\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__45723\,
            I => \N__45715\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__45720\,
            I => \N__45715\
        );

    \I__10711\ : Span4Mux_v
    port map (
            O => \N__45715\,
            I => \N__45710\
        );

    \I__10710\ : InMux
    port map (
            O => \N__45714\,
            I => \N__45707\
        );

    \I__10709\ : InMux
    port map (
            O => \N__45713\,
            I => \N__45704\
        );

    \I__10708\ : Span4Mux_h
    port map (
            O => \N__45710\,
            I => \N__45701\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__45707\,
            I => \N__45696\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__45704\,
            I => \N__45696\
        );

    \I__10705\ : Odrv4
    port map (
            O => \N__45701\,
            I => shift_flag_start
        );

    \I__10704\ : Odrv4
    port map (
            O => \N__45696\,
            I => shift_flag_start
        );

    \I__10703\ : IoInMux
    port map (
            O => \N__45691\,
            I => \N__45688\
        );

    \I__10702\ : LocalMux
    port map (
            O => \N__45688\,
            I => \N__45685\
        );

    \I__10701\ : Span4Mux_s1_v
    port map (
            O => \N__45685\,
            I => \N__45681\
        );

    \I__10700\ : InMux
    port map (
            O => \N__45684\,
            I => \N__45678\
        );

    \I__10699\ : Span4Mux_v
    port map (
            O => \N__45681\,
            I => \N__45673\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45673\
        );

    \I__10697\ : Span4Mux_v
    port map (
            O => \N__45673\,
            I => \N__45670\
        );

    \I__10696\ : Sp12to4
    port map (
            O => \N__45670\,
            I => \N__45667\
        );

    \I__10695\ : Span12Mux_h
    port map (
            O => \N__45667\,
            I => \N__45663\
        );

    \I__10694\ : InMux
    port map (
            O => \N__45666\,
            I => \N__45660\
        );

    \I__10693\ : Odrv12
    port map (
            O => \N__45663\,
            I => s3_phy_c
        );

    \I__10692\ : LocalMux
    port map (
            O => \N__45660\,
            I => s3_phy_c
        );

    \I__10691\ : CascadeMux
    port map (
            O => \N__45655\,
            I => \N__45644\
        );

    \I__10690\ : CascadeMux
    port map (
            O => \N__45654\,
            I => \N__45640\
        );

    \I__10689\ : CascadeMux
    port map (
            O => \N__45653\,
            I => \N__45637\
        );

    \I__10688\ : CascadeMux
    port map (
            O => \N__45652\,
            I => \N__45634\
        );

    \I__10687\ : CascadeMux
    port map (
            O => \N__45651\,
            I => \N__45631\
        );

    \I__10686\ : CascadeMux
    port map (
            O => \N__45650\,
            I => \N__45622\
        );

    \I__10685\ : CascadeMux
    port map (
            O => \N__45649\,
            I => \N__45615\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__45648\,
            I => \N__45612\
        );

    \I__10683\ : CascadeMux
    port map (
            O => \N__45647\,
            I => \N__45609\
        );

    \I__10682\ : InMux
    port map (
            O => \N__45644\,
            I => \N__45604\
        );

    \I__10681\ : InMux
    port map (
            O => \N__45643\,
            I => \N__45604\
        );

    \I__10680\ : InMux
    port map (
            O => \N__45640\,
            I => \N__45586\
        );

    \I__10679\ : InMux
    port map (
            O => \N__45637\,
            I => \N__45586\
        );

    \I__10678\ : InMux
    port map (
            O => \N__45634\,
            I => \N__45586\
        );

    \I__10677\ : InMux
    port map (
            O => \N__45631\,
            I => \N__45586\
        );

    \I__10676\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45586\
        );

    \I__10675\ : InMux
    port map (
            O => \N__45629\,
            I => \N__45586\
        );

    \I__10674\ : InMux
    port map (
            O => \N__45628\,
            I => \N__45586\
        );

    \I__10673\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45586\
        );

    \I__10672\ : InMux
    port map (
            O => \N__45626\,
            I => \N__45581\
        );

    \I__10671\ : InMux
    port map (
            O => \N__45625\,
            I => \N__45581\
        );

    \I__10670\ : InMux
    port map (
            O => \N__45622\,
            I => \N__45564\
        );

    \I__10669\ : InMux
    port map (
            O => \N__45621\,
            I => \N__45564\
        );

    \I__10668\ : InMux
    port map (
            O => \N__45620\,
            I => \N__45564\
        );

    \I__10667\ : InMux
    port map (
            O => \N__45619\,
            I => \N__45564\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45618\,
            I => \N__45564\
        );

    \I__10665\ : InMux
    port map (
            O => \N__45615\,
            I => \N__45564\
        );

    \I__10664\ : InMux
    port map (
            O => \N__45612\,
            I => \N__45564\
        );

    \I__10663\ : InMux
    port map (
            O => \N__45609\,
            I => \N__45564\
        );

    \I__10662\ : LocalMux
    port map (
            O => \N__45604\,
            I => \N__45561\
        );

    \I__10661\ : CascadeMux
    port map (
            O => \N__45603\,
            I => \N__45557\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__45586\,
            I => \N__45552\
        );

    \I__10659\ : LocalMux
    port map (
            O => \N__45581\,
            I => \N__45547\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__45564\,
            I => \N__45547\
        );

    \I__10657\ : Span4Mux_h
    port map (
            O => \N__45561\,
            I => \N__45544\
        );

    \I__10656\ : InMux
    port map (
            O => \N__45560\,
            I => \N__45541\
        );

    \I__10655\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45538\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45556\,
            I => \N__45533\
        );

    \I__10653\ : InMux
    port map (
            O => \N__45555\,
            I => \N__45533\
        );

    \I__10652\ : Span4Mux_h
    port map (
            O => \N__45552\,
            I => \N__45528\
        );

    \I__10651\ : Span4Mux_v
    port map (
            O => \N__45547\,
            I => \N__45528\
        );

    \I__10650\ : Span4Mux_h
    port map (
            O => \N__45544\,
            I => \N__45523\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__45541\,
            I => \N__45523\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__45538\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__45533\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10646\ : Odrv4
    port map (
            O => \N__45528\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10645\ : Odrv4
    port map (
            O => \N__45523\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__10644\ : InMux
    port map (
            O => \N__45514\,
            I => \N__45481\
        );

    \I__10643\ : InMux
    port map (
            O => \N__45513\,
            I => \N__45481\
        );

    \I__10642\ : InMux
    port map (
            O => \N__45512\,
            I => \N__45481\
        );

    \I__10641\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45481\
        );

    \I__10640\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45481\
        );

    \I__10639\ : InMux
    port map (
            O => \N__45509\,
            I => \N__45481\
        );

    \I__10638\ : InMux
    port map (
            O => \N__45508\,
            I => \N__45481\
        );

    \I__10637\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45481\
        );

    \I__10636\ : InMux
    port map (
            O => \N__45506\,
            I => \N__45464\
        );

    \I__10635\ : InMux
    port map (
            O => \N__45505\,
            I => \N__45464\
        );

    \I__10634\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45464\
        );

    \I__10633\ : InMux
    port map (
            O => \N__45503\,
            I => \N__45464\
        );

    \I__10632\ : InMux
    port map (
            O => \N__45502\,
            I => \N__45464\
        );

    \I__10631\ : InMux
    port map (
            O => \N__45501\,
            I => \N__45464\
        );

    \I__10630\ : InMux
    port map (
            O => \N__45500\,
            I => \N__45464\
        );

    \I__10629\ : InMux
    port map (
            O => \N__45499\,
            I => \N__45464\
        );

    \I__10628\ : CascadeMux
    port map (
            O => \N__45498\,
            I => \N__45461\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__45481\,
            I => \N__45451\
        );

    \I__10626\ : LocalMux
    port map (
            O => \N__45464\,
            I => \N__45451\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45446\
        );

    \I__10624\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45446\
        );

    \I__10623\ : InMux
    port map (
            O => \N__45459\,
            I => \N__45443\
        );

    \I__10622\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45438\
        );

    \I__10621\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45438\
        );

    \I__10620\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45435\
        );

    \I__10619\ : Span4Mux_v
    port map (
            O => \N__45451\,
            I => \N__45430\
        );

    \I__10618\ : LocalMux
    port map (
            O => \N__45446\,
            I => \N__45427\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__45443\,
            I => \N__45424\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__45438\,
            I => \N__45419\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__45435\,
            I => \N__45419\
        );

    \I__10614\ : InMux
    port map (
            O => \N__45434\,
            I => \N__45414\
        );

    \I__10613\ : InMux
    port map (
            O => \N__45433\,
            I => \N__45414\
        );

    \I__10612\ : Sp12to4
    port map (
            O => \N__45430\,
            I => \N__45409\
        );

    \I__10611\ : Span12Mux_v
    port map (
            O => \N__45427\,
            I => \N__45409\
        );

    \I__10610\ : Span4Mux_h
    port map (
            O => \N__45424\,
            I => \N__45406\
        );

    \I__10609\ : Span4Mux_h
    port map (
            O => \N__45419\,
            I => \N__45403\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__45414\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10607\ : Odrv12
    port map (
            O => \N__45409\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10606\ : Odrv4
    port map (
            O => \N__45406\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10605\ : Odrv4
    port map (
            O => \N__45403\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__10604\ : CascadeMux
    port map (
            O => \N__45394\,
            I => \N__45371\
        );

    \I__10603\ : InMux
    port map (
            O => \N__45393\,
            I => \N__45366\
        );

    \I__10602\ : InMux
    port map (
            O => \N__45392\,
            I => \N__45366\
        );

    \I__10601\ : CascadeMux
    port map (
            O => \N__45391\,
            I => \N__45362\
        );

    \I__10600\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45344\
        );

    \I__10599\ : InMux
    port map (
            O => \N__45389\,
            I => \N__45344\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45388\,
            I => \N__45344\
        );

    \I__10597\ : InMux
    port map (
            O => \N__45387\,
            I => \N__45344\
        );

    \I__10596\ : InMux
    port map (
            O => \N__45386\,
            I => \N__45344\
        );

    \I__10595\ : InMux
    port map (
            O => \N__45385\,
            I => \N__45344\
        );

    \I__10594\ : InMux
    port map (
            O => \N__45384\,
            I => \N__45344\
        );

    \I__10593\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45344\
        );

    \I__10592\ : InMux
    port map (
            O => \N__45382\,
            I => \N__45327\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45381\,
            I => \N__45327\
        );

    \I__10590\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45327\
        );

    \I__10589\ : InMux
    port map (
            O => \N__45379\,
            I => \N__45327\
        );

    \I__10588\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45327\
        );

    \I__10587\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45327\
        );

    \I__10586\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45327\
        );

    \I__10585\ : InMux
    port map (
            O => \N__45375\,
            I => \N__45327\
        );

    \I__10584\ : InMux
    port map (
            O => \N__45374\,
            I => \N__45323\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45371\,
            I => \N__45320\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__45366\,
            I => \N__45317\
        );

    \I__10581\ : InMux
    port map (
            O => \N__45365\,
            I => \N__45314\
        );

    \I__10580\ : InMux
    port map (
            O => \N__45362\,
            I => \N__45309\
        );

    \I__10579\ : InMux
    port map (
            O => \N__45361\,
            I => \N__45309\
        );

    \I__10578\ : LocalMux
    port map (
            O => \N__45344\,
            I => \N__45304\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__45327\,
            I => \N__45304\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45326\,
            I => \N__45301\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__45323\,
            I => \N__45292\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__45320\,
            I => \N__45292\
        );

    \I__10573\ : Span4Mux_v
    port map (
            O => \N__45317\,
            I => \N__45292\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__45314\,
            I => \N__45292\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__45309\,
            I => \N__45287\
        );

    \I__10570\ : Span4Mux_v
    port map (
            O => \N__45304\,
            I => \N__45287\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__45301\,
            I => \N__45284\
        );

    \I__10568\ : Span4Mux_h
    port map (
            O => \N__45292\,
            I => \N__45281\
        );

    \I__10567\ : Odrv4
    port map (
            O => \N__45287\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10566\ : Odrv12
    port map (
            O => \N__45284\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10565\ : Odrv4
    port map (
            O => \N__45281\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__10564\ : InMux
    port map (
            O => \N__45274\,
            I => \N__45271\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__45271\,
            I => \N__45267\
        );

    \I__10562\ : InMux
    port map (
            O => \N__45270\,
            I => \N__45264\
        );

    \I__10561\ : Span4Mux_h
    port map (
            O => \N__45267\,
            I => \N__45260\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__45264\,
            I => \N__45257\
        );

    \I__10559\ : InMux
    port map (
            O => \N__45263\,
            I => \N__45254\
        );

    \I__10558\ : Span4Mux_v
    port map (
            O => \N__45260\,
            I => \N__45250\
        );

    \I__10557\ : Span12Mux_s11_v
    port map (
            O => \N__45257\,
            I => \N__45245\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__45254\,
            I => \N__45245\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45253\,
            I => \N__45242\
        );

    \I__10554\ : Odrv4
    port map (
            O => \N__45250\,
            I => measured_delay_tr_16
        );

    \I__10553\ : Odrv12
    port map (
            O => \N__45245\,
            I => measured_delay_tr_16
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__45242\,
            I => measured_delay_tr_16
        );

    \I__10551\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45232\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__45232\,
            I => \N__45229\
        );

    \I__10549\ : Span4Mux_h
    port map (
            O => \N__45229\,
            I => \N__45226\
        );

    \I__10548\ : Odrv4
    port map (
            O => \N__45226\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__10547\ : CEMux
    port map (
            O => \N__45223\,
            I => \N__45220\
        );

    \I__10546\ : LocalMux
    port map (
            O => \N__45220\,
            I => \N__45216\
        );

    \I__10545\ : CEMux
    port map (
            O => \N__45219\,
            I => \N__45213\
        );

    \I__10544\ : Span4Mux_v
    port map (
            O => \N__45216\,
            I => \N__45206\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__45213\,
            I => \N__45206\
        );

    \I__10542\ : CEMux
    port map (
            O => \N__45212\,
            I => \N__45203\
        );

    \I__10541\ : CEMux
    port map (
            O => \N__45211\,
            I => \N__45200\
        );

    \I__10540\ : Span4Mux_h
    port map (
            O => \N__45206\,
            I => \N__45197\
        );

    \I__10539\ : LocalMux
    port map (
            O => \N__45203\,
            I => \N__45193\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__45200\,
            I => \N__45190\
        );

    \I__10537\ : Span4Mux_h
    port map (
            O => \N__45197\,
            I => \N__45187\
        );

    \I__10536\ : CEMux
    port map (
            O => \N__45196\,
            I => \N__45184\
        );

    \I__10535\ : Span4Mux_h
    port map (
            O => \N__45193\,
            I => \N__45181\
        );

    \I__10534\ : Span4Mux_h
    port map (
            O => \N__45190\,
            I => \N__45176\
        );

    \I__10533\ : Span4Mux_v
    port map (
            O => \N__45187\,
            I => \N__45176\
        );

    \I__10532\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45173\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__45181\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__45176\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10529\ : Odrv12
    port map (
            O => \N__45173\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__45166\,
            I => \N__45161\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__45165\,
            I => \N__45158\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45164\,
            I => \N__45142\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45161\,
            I => \N__45142\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45158\,
            I => \N__45142\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45157\,
            I => \N__45142\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45156\,
            I => \N__45142\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45138\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45154\,
            I => \N__45128\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45153\,
            I => \N__45125\
        );

    \I__10518\ : LocalMux
    port map (
            O => \N__45142\,
            I => \N__45122\
        );

    \I__10517\ : InMux
    port map (
            O => \N__45141\,
            I => \N__45119\
        );

    \I__10516\ : LocalMux
    port map (
            O => \N__45138\,
            I => \N__45116\
        );

    \I__10515\ : InMux
    port map (
            O => \N__45137\,
            I => \N__45113\
        );

    \I__10514\ : InMux
    port map (
            O => \N__45136\,
            I => \N__45106\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45106\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45106\
        );

    \I__10511\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45099\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45099\
        );

    \I__10509\ : InMux
    port map (
            O => \N__45131\,
            I => \N__45099\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45128\,
            I => \N__45094\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__45125\,
            I => \N__45094\
        );

    \I__10506\ : Span4Mux_h
    port map (
            O => \N__45122\,
            I => \N__45089\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__45119\,
            I => \N__45089\
        );

    \I__10504\ : Span4Mux_v
    port map (
            O => \N__45116\,
            I => \N__45084\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45084\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__45106\,
            I => \N__45079\
        );

    \I__10501\ : LocalMux
    port map (
            O => \N__45099\,
            I => \N__45079\
        );

    \I__10500\ : Span4Mux_h
    port map (
            O => \N__45094\,
            I => \N__45076\
        );

    \I__10499\ : Span4Mux_v
    port map (
            O => \N__45089\,
            I => \N__45071\
        );

    \I__10498\ : Span4Mux_h
    port map (
            O => \N__45084\,
            I => \N__45071\
        );

    \I__10497\ : Span4Mux_h
    port map (
            O => \N__45079\,
            I => \N__45068\
        );

    \I__10496\ : Span4Mux_h
    port map (
            O => \N__45076\,
            I => \N__45065\
        );

    \I__10495\ : Odrv4
    port map (
            O => \N__45071\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__10494\ : Odrv4
    port map (
            O => \N__45068\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__10493\ : Odrv4
    port map (
            O => \N__45065\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__10492\ : CascadeMux
    port map (
            O => \N__45058\,
            I => \N__45054\
        );

    \I__10491\ : InMux
    port map (
            O => \N__45057\,
            I => \N__45049\
        );

    \I__10490\ : InMux
    port map (
            O => \N__45054\,
            I => \N__45044\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45053\,
            I => \N__45044\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45052\,
            I => \N__45041\
        );

    \I__10487\ : LocalMux
    port map (
            O => \N__45049\,
            I => \N__45038\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__45044\,
            I => \N__45035\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45041\,
            I => \N__45030\
        );

    \I__10484\ : Span4Mux_v
    port map (
            O => \N__45038\,
            I => \N__45027\
        );

    \I__10483\ : Span12Mux_h
    port map (
            O => \N__45035\,
            I => \N__45024\
        );

    \I__10482\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45019\
        );

    \I__10481\ : InMux
    port map (
            O => \N__45033\,
            I => \N__45019\
        );

    \I__10480\ : Span4Mux_h
    port map (
            O => \N__45030\,
            I => \N__45014\
        );

    \I__10479\ : Span4Mux_h
    port map (
            O => \N__45027\,
            I => \N__45014\
        );

    \I__10478\ : Odrv12
    port map (
            O => \N__45024\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45019\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__10476\ : Odrv4
    port map (
            O => \N__45014\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45007\,
            I => \N__44995\
        );

    \I__10474\ : InMux
    port map (
            O => \N__45006\,
            I => \N__44995\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45005\,
            I => \N__44995\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45004\,
            I => \N__44995\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__44995\,
            I => \N__44990\
        );

    \I__10470\ : InMux
    port map (
            O => \N__44994\,
            I => \N__44987\
        );

    \I__10469\ : InMux
    port map (
            O => \N__44993\,
            I => \N__44984\
        );

    \I__10468\ : Span4Mux_h
    port map (
            O => \N__44990\,
            I => \N__44979\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__44987\,
            I => \N__44979\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__44984\,
            I => \N__44976\
        );

    \I__10465\ : Span4Mux_v
    port map (
            O => \N__44979\,
            I => \N__44969\
        );

    \I__10464\ : Span4Mux_v
    port map (
            O => \N__44976\,
            I => \N__44966\
        );

    \I__10463\ : InMux
    port map (
            O => \N__44975\,
            I => \N__44963\
        );

    \I__10462\ : InMux
    port map (
            O => \N__44974\,
            I => \N__44956\
        );

    \I__10461\ : InMux
    port map (
            O => \N__44973\,
            I => \N__44956\
        );

    \I__10460\ : InMux
    port map (
            O => \N__44972\,
            I => \N__44956\
        );

    \I__10459\ : Span4Mux_h
    port map (
            O => \N__44969\,
            I => \N__44953\
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__44966\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__10457\ : LocalMux
    port map (
            O => \N__44963\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__10456\ : LocalMux
    port map (
            O => \N__44956\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__44953\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\
        );

    \I__10454\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44940\
        );

    \I__10453\ : InMux
    port map (
            O => \N__44943\,
            I => \N__44937\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__44940\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__44937\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10450\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44929\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__44929\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__10448\ : InMux
    port map (
            O => \N__44926\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__10447\ : InMux
    port map (
            O => \N__44923\,
            I => \N__44919\
        );

    \I__10446\ : InMux
    port map (
            O => \N__44922\,
            I => \N__44916\
        );

    \I__10445\ : LocalMux
    port map (
            O => \N__44919\,
            I => \N__44913\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__44916\,
            I => \N__44910\
        );

    \I__10443\ : Odrv4
    port map (
            O => \N__44913\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10442\ : Odrv4
    port map (
            O => \N__44910\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10441\ : CascadeMux
    port map (
            O => \N__44905\,
            I => \N__44902\
        );

    \I__10440\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44899\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__44899\,
            I => \N__44896\
        );

    \I__10438\ : Odrv4
    port map (
            O => \N__44896\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__10437\ : InMux
    port map (
            O => \N__44893\,
            I => \bfn_18_10_0_\
        );

    \I__10436\ : InMux
    port map (
            O => \N__44890\,
            I => \N__44886\
        );

    \I__10435\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44883\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__44886\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__44883\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__10432\ : InMux
    port map (
            O => \N__44878\,
            I => \N__44875\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__44875\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__10430\ : InMux
    port map (
            O => \N__44872\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__10429\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44866\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__44866\,
            I => \N__44862\
        );

    \I__10427\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44859\
        );

    \I__10426\ : Span4Mux_h
    port map (
            O => \N__44862\,
            I => \N__44854\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__44859\,
            I => \N__44854\
        );

    \I__10424\ : Span4Mux_h
    port map (
            O => \N__44854\,
            I => \N__44851\
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__44851\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__10422\ : InMux
    port map (
            O => \N__44848\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__10421\ : InMux
    port map (
            O => \N__44845\,
            I => \N__44842\
        );

    \I__10420\ : LocalMux
    port map (
            O => \N__44842\,
            I => \N__44839\
        );

    \I__10419\ : Span4Mux_v
    port map (
            O => \N__44839\,
            I => \N__44836\
        );

    \I__10418\ : Odrv4
    port map (
            O => \N__44836\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__10417\ : InMux
    port map (
            O => \N__44833\,
            I => \N__44830\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__44830\,
            I => \N__44827\
        );

    \I__10415\ : Odrv4
    port map (
            O => \N__44827\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa\
        );

    \I__10414\ : InMux
    port map (
            O => \N__44824\,
            I => \N__44818\
        );

    \I__10413\ : InMux
    port map (
            O => \N__44823\,
            I => \N__44811\
        );

    \I__10412\ : InMux
    port map (
            O => \N__44822\,
            I => \N__44811\
        );

    \I__10411\ : InMux
    port map (
            O => \N__44821\,
            I => \N__44811\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__44818\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__10409\ : LocalMux
    port map (
            O => \N__44811\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__10408\ : CascadeMux
    port map (
            O => \N__44806\,
            I => \N__44802\
        );

    \I__10407\ : CascadeMux
    port map (
            O => \N__44805\,
            I => \N__44799\
        );

    \I__10406\ : InMux
    port map (
            O => \N__44802\,
            I => \N__44795\
        );

    \I__10405\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44790\
        );

    \I__10404\ : InMux
    port map (
            O => \N__44798\,
            I => \N__44790\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__44795\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__10402\ : LocalMux
    port map (
            O => \N__44790\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__10401\ : IoInMux
    port map (
            O => \N__44785\,
            I => \N__44782\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__44782\,
            I => \N__44779\
        );

    \I__10399\ : IoSpan4Mux
    port map (
            O => \N__44779\,
            I => \N__44776\
        );

    \I__10398\ : Span4Mux_s3_v
    port map (
            O => \N__44776\,
            I => \N__44773\
        );

    \I__10397\ : Span4Mux_v
    port map (
            O => \N__44773\,
            I => \N__44770\
        );

    \I__10396\ : Sp12to4
    port map (
            O => \N__44770\,
            I => \N__44767\
        );

    \I__10395\ : Span12Mux_h
    port map (
            O => \N__44767\,
            I => \N__44763\
        );

    \I__10394\ : CascadeMux
    port map (
            O => \N__44766\,
            I => \N__44760\
        );

    \I__10393\ : Span12Mux_v
    port map (
            O => \N__44763\,
            I => \N__44757\
        );

    \I__10392\ : InMux
    port map (
            O => \N__44760\,
            I => \N__44754\
        );

    \I__10391\ : Odrv12
    port map (
            O => \N__44757\,
            I => s4_phy_c
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__44754\,
            I => s4_phy_c
        );

    \I__10389\ : InMux
    port map (
            O => \N__44749\,
            I => \N__44745\
        );

    \I__10388\ : InMux
    port map (
            O => \N__44748\,
            I => \N__44742\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__44745\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10386\ : LocalMux
    port map (
            O => \N__44742\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__10385\ : InMux
    port map (
            O => \N__44737\,
            I => \N__44734\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__44734\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__10383\ : InMux
    port map (
            O => \N__44731\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__10382\ : InMux
    port map (
            O => \N__44728\,
            I => \N__44725\
        );

    \I__10381\ : LocalMux
    port map (
            O => \N__44725\,
            I => \N__44722\
        );

    \I__10380\ : Span4Mux_h
    port map (
            O => \N__44722\,
            I => \N__44718\
        );

    \I__10379\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44715\
        );

    \I__10378\ : Odrv4
    port map (
            O => \N__44718\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__44715\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__10376\ : InMux
    port map (
            O => \N__44710\,
            I => \N__44707\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44704\
        );

    \I__10374\ : Span4Mux_h
    port map (
            O => \N__44704\,
            I => \N__44701\
        );

    \I__10373\ : Odrv4
    port map (
            O => \N__44701\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__10372\ : InMux
    port map (
            O => \N__44698\,
            I => \bfn_18_9_0_\
        );

    \I__10371\ : InMux
    port map (
            O => \N__44695\,
            I => \N__44691\
        );

    \I__10370\ : InMux
    port map (
            O => \N__44694\,
            I => \N__44688\
        );

    \I__10369\ : LocalMux
    port map (
            O => \N__44691\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__44688\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__10367\ : InMux
    port map (
            O => \N__44683\,
            I => \N__44680\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__44680\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44677\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__10364\ : InMux
    port map (
            O => \N__44674\,
            I => \N__44670\
        );

    \I__10363\ : InMux
    port map (
            O => \N__44673\,
            I => \N__44667\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44670\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__44667\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__10360\ : InMux
    port map (
            O => \N__44662\,
            I => \N__44659\
        );

    \I__10359\ : LocalMux
    port map (
            O => \N__44659\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__10358\ : InMux
    port map (
            O => \N__44656\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__10357\ : InMux
    port map (
            O => \N__44653\,
            I => \N__44649\
        );

    \I__10356\ : InMux
    port map (
            O => \N__44652\,
            I => \N__44646\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__44649\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10354\ : LocalMux
    port map (
            O => \N__44646\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__10353\ : InMux
    port map (
            O => \N__44641\,
            I => \N__44638\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__44638\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__10351\ : InMux
    port map (
            O => \N__44635\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__10350\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44628\
        );

    \I__10349\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44625\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__44628\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10347\ : LocalMux
    port map (
            O => \N__44625\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__10346\ : InMux
    port map (
            O => \N__44620\,
            I => \N__44617\
        );

    \I__10345\ : LocalMux
    port map (
            O => \N__44617\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__10344\ : InMux
    port map (
            O => \N__44614\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__10343\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44607\
        );

    \I__10342\ : InMux
    port map (
            O => \N__44610\,
            I => \N__44604\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__44607\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__44604\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__10339\ : InMux
    port map (
            O => \N__44599\,
            I => \N__44596\
        );

    \I__10338\ : LocalMux
    port map (
            O => \N__44596\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__10337\ : InMux
    port map (
            O => \N__44593\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__10336\ : InMux
    port map (
            O => \N__44590\,
            I => \N__44586\
        );

    \I__10335\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44583\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__44586\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__44583\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__10332\ : InMux
    port map (
            O => \N__44578\,
            I => \N__44575\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__44575\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__10330\ : InMux
    port map (
            O => \N__44572\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__10329\ : InMux
    port map (
            O => \N__44569\,
            I => \N__44531\
        );

    \I__10328\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44531\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44567\,
            I => \N__44531\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44566\,
            I => \N__44531\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44565\,
            I => \N__44526\
        );

    \I__10324\ : InMux
    port map (
            O => \N__44564\,
            I => \N__44526\
        );

    \I__10323\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44517\
        );

    \I__10322\ : InMux
    port map (
            O => \N__44562\,
            I => \N__44517\
        );

    \I__10321\ : InMux
    port map (
            O => \N__44561\,
            I => \N__44517\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44560\,
            I => \N__44517\
        );

    \I__10319\ : InMux
    port map (
            O => \N__44559\,
            I => \N__44508\
        );

    \I__10318\ : InMux
    port map (
            O => \N__44558\,
            I => \N__44508\
        );

    \I__10317\ : InMux
    port map (
            O => \N__44557\,
            I => \N__44508\
        );

    \I__10316\ : InMux
    port map (
            O => \N__44556\,
            I => \N__44508\
        );

    \I__10315\ : InMux
    port map (
            O => \N__44555\,
            I => \N__44499\
        );

    \I__10314\ : InMux
    port map (
            O => \N__44554\,
            I => \N__44499\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44499\
        );

    \I__10312\ : InMux
    port map (
            O => \N__44552\,
            I => \N__44499\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44551\,
            I => \N__44490\
        );

    \I__10310\ : InMux
    port map (
            O => \N__44550\,
            I => \N__44490\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44549\,
            I => \N__44490\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44490\
        );

    \I__10307\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44481\
        );

    \I__10306\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44481\
        );

    \I__10305\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44481\
        );

    \I__10304\ : InMux
    port map (
            O => \N__44544\,
            I => \N__44481\
        );

    \I__10303\ : InMux
    port map (
            O => \N__44543\,
            I => \N__44472\
        );

    \I__10302\ : InMux
    port map (
            O => \N__44542\,
            I => \N__44472\
        );

    \I__10301\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44472\
        );

    \I__10300\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44472\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__44531\,
            I => \N__44461\
        );

    \I__10298\ : LocalMux
    port map (
            O => \N__44526\,
            I => \N__44461\
        );

    \I__10297\ : LocalMux
    port map (
            O => \N__44517\,
            I => \N__44461\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__44508\,
            I => \N__44461\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__44499\,
            I => \N__44461\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__44490\,
            I => \N__44458\
        );

    \I__10293\ : LocalMux
    port map (
            O => \N__44481\,
            I => \N__44451\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__44472\,
            I => \N__44451\
        );

    \I__10291\ : Span4Mux_v
    port map (
            O => \N__44461\,
            I => \N__44451\
        );

    \I__10290\ : Odrv12
    port map (
            O => \N__44458\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__10289\ : Odrv4
    port map (
            O => \N__44451\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__10288\ : InMux
    port map (
            O => \N__44446\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__10287\ : CEMux
    port map (
            O => \N__44443\,
            I => \N__44437\
        );

    \I__10286\ : CEMux
    port map (
            O => \N__44442\,
            I => \N__44434\
        );

    \I__10285\ : CEMux
    port map (
            O => \N__44441\,
            I => \N__44431\
        );

    \I__10284\ : CEMux
    port map (
            O => \N__44440\,
            I => \N__44428\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__44437\,
            I => \N__44425\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__44434\,
            I => \N__44422\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__44431\,
            I => \N__44417\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__44428\,
            I => \N__44417\
        );

    \I__10279\ : Span4Mux_v
    port map (
            O => \N__44425\,
            I => \N__44410\
        );

    \I__10278\ : Span4Mux_v
    port map (
            O => \N__44422\,
            I => \N__44410\
        );

    \I__10277\ : Span4Mux_v
    port map (
            O => \N__44417\,
            I => \N__44410\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__44410\,
            I => \delay_measurement_inst.delay_tr_timer.N_339_i\
        );

    \I__10275\ : InMux
    port map (
            O => \N__44407\,
            I => \N__44404\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__44404\,
            I => \N__44401\
        );

    \I__10273\ : Odrv4
    port map (
            O => \N__44401\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__10272\ : CascadeMux
    port map (
            O => \N__44398\,
            I => \N__44394\
        );

    \I__10271\ : InMux
    port map (
            O => \N__44397\,
            I => \N__44390\
        );

    \I__10270\ : InMux
    port map (
            O => \N__44394\,
            I => \N__44387\
        );

    \I__10269\ : InMux
    port map (
            O => \N__44393\,
            I => \N__44384\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__44390\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10267\ : LocalMux
    port map (
            O => \N__44387\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10266\ : LocalMux
    port map (
            O => \N__44384\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__10265\ : InMux
    port map (
            O => \N__44377\,
            I => \N__44373\
        );

    \I__10264\ : InMux
    port map (
            O => \N__44376\,
            I => \N__44370\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__44373\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10262\ : LocalMux
    port map (
            O => \N__44370\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__10261\ : InMux
    port map (
            O => \N__44365\,
            I => \N__44362\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__44362\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__10259\ : InMux
    port map (
            O => \N__44359\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__10258\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44353\
        );

    \I__10257\ : LocalMux
    port map (
            O => \N__44353\,
            I => \N__44350\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__44350\,
            I => \N__44347\
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__44347\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\
        );

    \I__10254\ : CascadeMux
    port map (
            O => \N__44344\,
            I => \N__44341\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44341\,
            I => \N__44337\
        );

    \I__10252\ : InMux
    port map (
            O => \N__44340\,
            I => \N__44334\
        );

    \I__10251\ : LocalMux
    port map (
            O => \N__44337\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__44334\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__10249\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44326\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__44326\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__10247\ : InMux
    port map (
            O => \N__44323\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__10246\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44316\
        );

    \I__10245\ : InMux
    port map (
            O => \N__44319\,
            I => \N__44313\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__44316\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__44313\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__10242\ : CascadeMux
    port map (
            O => \N__44308\,
            I => \N__44305\
        );

    \I__10241\ : InMux
    port map (
            O => \N__44305\,
            I => \N__44302\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__44302\,
            I => \N__44299\
        );

    \I__10239\ : Odrv4
    port map (
            O => \N__44299\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44296\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44293\,
            I => \N__44289\
        );

    \I__10236\ : InMux
    port map (
            O => \N__44292\,
            I => \N__44286\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__44289\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__44286\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__10233\ : CascadeMux
    port map (
            O => \N__44281\,
            I => \N__44278\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44278\,
            I => \N__44275\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__44275\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44272\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44269\,
            I => \N__44265\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44268\,
            I => \N__44262\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__44265\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10226\ : LocalMux
    port map (
            O => \N__44262\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44257\,
            I => \N__44254\
        );

    \I__10224\ : LocalMux
    port map (
            O => \N__44254\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44251\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44248\,
            I => \N__44245\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__44245\,
            I => \N__44241\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44238\
        );

    \I__10219\ : Span4Mux_h
    port map (
            O => \N__44241\,
            I => \N__44235\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__44238\,
            I => \N__44232\
        );

    \I__10217\ : Odrv4
    port map (
            O => \N__44235\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10216\ : Odrv4
    port map (
            O => \N__44232\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44227\,
            I => \N__44224\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__44224\,
            I => \N__44221\
        );

    \I__10213\ : Span4Mux_h
    port map (
            O => \N__44221\,
            I => \N__44218\
        );

    \I__10212\ : Odrv4
    port map (
            O => \N__44218\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__10211\ : InMux
    port map (
            O => \N__44215\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__10210\ : InMux
    port map (
            O => \N__44212\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__10209\ : InMux
    port map (
            O => \N__44209\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__10208\ : InMux
    port map (
            O => \N__44206\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44203\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44200\,
            I => \bfn_17_26_0_\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44197\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__10204\ : InMux
    port map (
            O => \N__44194\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__10203\ : InMux
    port map (
            O => \N__44191\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__10202\ : InMux
    port map (
            O => \N__44188\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44185\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__10200\ : InMux
    port map (
            O => \N__44182\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44179\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44176\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__10197\ : InMux
    port map (
            O => \N__44173\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44170\,
            I => \bfn_17_25_0_\
        );

    \I__10195\ : InMux
    port map (
            O => \N__44167\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44164\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44161\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44158\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44155\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44152\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44149\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44146\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44143\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44140\,
            I => \bfn_17_24_0_\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44137\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44134\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44131\,
            I => \N__44128\
        );

    \I__10182\ : LocalMux
    port map (
            O => \N__44128\,
            I => \N__44124\
        );

    \I__10181\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44121\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__44124\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10179\ : LocalMux
    port map (
            O => \N__44121\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44116\,
            I => \N__44111\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44115\,
            I => \N__44108\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44114\,
            I => \N__44105\
        );

    \I__10175\ : LocalMux
    port map (
            O => \N__44111\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44108\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44105\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44098\,
            I => \N__44094\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44097\,
            I => \N__44091\
        );

    \I__10170\ : LocalMux
    port map (
            O => \N__44094\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\
        );

    \I__10169\ : LocalMux
    port map (
            O => \N__44091\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\
        );

    \I__10168\ : CascadeMux
    port map (
            O => \N__44086\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44083\,
            I => \N__44068\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44082\,
            I => \N__44068\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44081\,
            I => \N__44068\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44080\,
            I => \N__44068\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44079\,
            I => \N__44068\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44068\,
            I => \N__44065\
        );

    \I__10161\ : Span4Mux_h
    port map (
            O => \N__44065\,
            I => \N__44062\
        );

    \I__10160\ : Odrv4
    port map (
            O => \N__44062\,
            I => \delay_measurement_inst.N_409_1\
        );

    \I__10159\ : InMux
    port map (
            O => \N__44059\,
            I => \N__44053\
        );

    \I__10158\ : InMux
    port map (
            O => \N__44058\,
            I => \N__44050\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44057\,
            I => \N__44045\
        );

    \I__10156\ : InMux
    port map (
            O => \N__44056\,
            I => \N__44045\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44053\,
            I => \N__44042\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44050\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__10153\ : LocalMux
    port map (
            O => \N__44045\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__10152\ : Odrv4
    port map (
            O => \N__44042\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__10151\ : CascadeMux
    port map (
            O => \N__44035\,
            I => \N__44032\
        );

    \I__10150\ : InMux
    port map (
            O => \N__44032\,
            I => \N__44029\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__44029\,
            I => \N__44026\
        );

    \I__10148\ : Span4Mux_h
    port map (
            O => \N__44026\,
            I => \N__44023\
        );

    \I__10147\ : Odrv4
    port map (
            O => \N__44023\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44020\,
            I => \bfn_17_23_0_\
        );

    \I__10145\ : InMux
    port map (
            O => \N__44017\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44011\
        );

    \I__10143\ : LocalMux
    port map (
            O => \N__44011\,
            I => \N__44007\
        );

    \I__10142\ : InMux
    port map (
            O => \N__44010\,
            I => \N__44003\
        );

    \I__10141\ : Span4Mux_v
    port map (
            O => \N__44007\,
            I => \N__44000\
        );

    \I__10140\ : InMux
    port map (
            O => \N__44006\,
            I => \N__43997\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__44003\,
            I => \N__43994\
        );

    \I__10138\ : Odrv4
    port map (
            O => \N__44000\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__43997\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__10136\ : Odrv12
    port map (
            O => \N__43994\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__10135\ : InMux
    port map (
            O => \N__43987\,
            I => \N__43982\
        );

    \I__10134\ : InMux
    port map (
            O => \N__43986\,
            I => \N__43976\
        );

    \I__10133\ : InMux
    port map (
            O => \N__43985\,
            I => \N__43976\
        );

    \I__10132\ : LocalMux
    port map (
            O => \N__43982\,
            I => \N__43973\
        );

    \I__10131\ : InMux
    port map (
            O => \N__43981\,
            I => \N__43970\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__43976\,
            I => \N__43967\
        );

    \I__10129\ : Sp12to4
    port map (
            O => \N__43973\,
            I => \N__43962\
        );

    \I__10128\ : LocalMux
    port map (
            O => \N__43970\,
            I => \N__43962\
        );

    \I__10127\ : Span12Mux_v
    port map (
            O => \N__43967\,
            I => \N__43959\
        );

    \I__10126\ : Span12Mux_v
    port map (
            O => \N__43962\,
            I => \N__43956\
        );

    \I__10125\ : Odrv12
    port map (
            O => \N__43959\,
            I => delay_tr_d2
        );

    \I__10124\ : Odrv12
    port map (
            O => \N__43956\,
            I => delay_tr_d2
        );

    \I__10123\ : InMux
    port map (
            O => \N__43951\,
            I => \N__43948\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43944\
        );

    \I__10121\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43940\
        );

    \I__10120\ : Span4Mux_h
    port map (
            O => \N__43944\,
            I => \N__43937\
        );

    \I__10119\ : InMux
    port map (
            O => \N__43943\,
            I => \N__43934\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__43940\,
            I => \N__43931\
        );

    \I__10117\ : Odrv4
    port map (
            O => \N__43937\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__43934\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__10115\ : Odrv12
    port map (
            O => \N__43931\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__10114\ : CascadeMux
    port map (
            O => \N__43924\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4_cascade_\
        );

    \I__10113\ : InMux
    port map (
            O => \N__43921\,
            I => \N__43918\
        );

    \I__10112\ : LocalMux
    port map (
            O => \N__43918\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5\
        );

    \I__10111\ : CascadeMux
    port map (
            O => \N__43915\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\
        );

    \I__10110\ : InMux
    port map (
            O => \N__43912\,
            I => \N__43909\
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__43909\,
            I => \N__43905\
        );

    \I__10108\ : InMux
    port map (
            O => \N__43908\,
            I => \N__43902\
        );

    \I__10107\ : Span4Mux_h
    port map (
            O => \N__43905\,
            I => \N__43899\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__43902\,
            I => \N__43896\
        );

    \I__10105\ : Span4Mux_h
    port map (
            O => \N__43899\,
            I => \N__43893\
        );

    \I__10104\ : Odrv12
    port map (
            O => \N__43896\,
            I => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\
        );

    \I__10103\ : Odrv4
    port map (
            O => \N__43893\,
            I => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\
        );

    \I__10102\ : CascadeMux
    port map (
            O => \N__43888\,
            I => \delay_measurement_inst.delay_tr_timer.N_390_cascade_\
        );

    \I__10101\ : InMux
    port map (
            O => \N__43885\,
            I => \N__43882\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__43882\,
            I => \delay_measurement_inst.delay_tr_timer.N_379\
        );

    \I__10099\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43873\
        );

    \I__10098\ : InMux
    port map (
            O => \N__43878\,
            I => \N__43870\
        );

    \I__10097\ : InMux
    port map (
            O => \N__43877\,
            I => \N__43865\
        );

    \I__10096\ : InMux
    port map (
            O => \N__43876\,
            I => \N__43865\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__43873\,
            I => \N__43860\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__43870\,
            I => \N__43860\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__43865\,
            I => \N__43857\
        );

    \I__10092\ : Span4Mux_v
    port map (
            O => \N__43860\,
            I => \N__43852\
        );

    \I__10091\ : Span4Mux_v
    port map (
            O => \N__43857\,
            I => \N__43852\
        );

    \I__10090\ : Span4Mux_h
    port map (
            O => \N__43852\,
            I => \N__43848\
        );

    \I__10089\ : InMux
    port map (
            O => \N__43851\,
            I => \N__43845\
        );

    \I__10088\ : Odrv4
    port map (
            O => \N__43848\,
            I => \delay_measurement_inst.N_280_i\
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__43845\,
            I => \delay_measurement_inst.N_280_i\
        );

    \I__10086\ : InMux
    port map (
            O => \N__43840\,
            I => \bfn_17_14_0_\
        );

    \I__10085\ : CascadeMux
    port map (
            O => \N__43837\,
            I => \N__43833\
        );

    \I__10084\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43830\
        );

    \I__10083\ : InMux
    port map (
            O => \N__43833\,
            I => \N__43827\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__43830\,
            I => \N__43821\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__43827\,
            I => \N__43821\
        );

    \I__10080\ : InMux
    port map (
            O => \N__43826\,
            I => \N__43818\
        );

    \I__10079\ : Span4Mux_v
    port map (
            O => \N__43821\,
            I => \N__43815\
        );

    \I__10078\ : LocalMux
    port map (
            O => \N__43818\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10077\ : Odrv4
    port map (
            O => \N__43815\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10076\ : InMux
    port map (
            O => \N__43810\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__10075\ : CascadeMux
    port map (
            O => \N__43807\,
            I => \N__43803\
        );

    \I__10074\ : CascadeMux
    port map (
            O => \N__43806\,
            I => \N__43800\
        );

    \I__10073\ : InMux
    port map (
            O => \N__43803\,
            I => \N__43794\
        );

    \I__10072\ : InMux
    port map (
            O => \N__43800\,
            I => \N__43794\
        );

    \I__10071\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43791\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__43794\,
            I => \N__43788\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__43791\,
            I => \N__43783\
        );

    \I__10068\ : Span4Mux_v
    port map (
            O => \N__43788\,
            I => \N__43783\
        );

    \I__10067\ : Odrv4
    port map (
            O => \N__43783\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__10066\ : InMux
    port map (
            O => \N__43780\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__10065\ : CascadeMux
    port map (
            O => \N__43777\,
            I => \N__43773\
        );

    \I__10064\ : InMux
    port map (
            O => \N__43776\,
            I => \N__43769\
        );

    \I__10063\ : InMux
    port map (
            O => \N__43773\,
            I => \N__43766\
        );

    \I__10062\ : InMux
    port map (
            O => \N__43772\,
            I => \N__43763\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__43769\,
            I => \N__43758\
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__43766\,
            I => \N__43758\
        );

    \I__10059\ : LocalMux
    port map (
            O => \N__43763\,
            I => \N__43753\
        );

    \I__10058\ : Span4Mux_v
    port map (
            O => \N__43758\,
            I => \N__43753\
        );

    \I__10057\ : Odrv4
    port map (
            O => \N__43753\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10056\ : InMux
    port map (
            O => \N__43750\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__10055\ : InMux
    port map (
            O => \N__43747\,
            I => \N__43744\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__43744\,
            I => \N__43740\
        );

    \I__10053\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43737\
        );

    \I__10052\ : Span4Mux_v
    port map (
            O => \N__43740\,
            I => \N__43734\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__43737\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10050\ : Odrv4
    port map (
            O => \N__43734\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10049\ : InMux
    port map (
            O => \N__43729\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43726\,
            I => \N__43694\
        );

    \I__10047\ : InMux
    port map (
            O => \N__43725\,
            I => \N__43694\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43724\,
            I => \N__43694\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43723\,
            I => \N__43694\
        );

    \I__10044\ : InMux
    port map (
            O => \N__43722\,
            I => \N__43685\
        );

    \I__10043\ : InMux
    port map (
            O => \N__43721\,
            I => \N__43685\
        );

    \I__10042\ : InMux
    port map (
            O => \N__43720\,
            I => \N__43685\
        );

    \I__10041\ : InMux
    port map (
            O => \N__43719\,
            I => \N__43685\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43718\,
            I => \N__43676\
        );

    \I__10039\ : InMux
    port map (
            O => \N__43717\,
            I => \N__43676\
        );

    \I__10038\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43676\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43715\,
            I => \N__43676\
        );

    \I__10036\ : InMux
    port map (
            O => \N__43714\,
            I => \N__43667\
        );

    \I__10035\ : InMux
    port map (
            O => \N__43713\,
            I => \N__43667\
        );

    \I__10034\ : InMux
    port map (
            O => \N__43712\,
            I => \N__43667\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43711\,
            I => \N__43667\
        );

    \I__10032\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43658\
        );

    \I__10031\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43658\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43708\,
            I => \N__43658\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43707\,
            I => \N__43658\
        );

    \I__10028\ : InMux
    port map (
            O => \N__43706\,
            I => \N__43649\
        );

    \I__10027\ : InMux
    port map (
            O => \N__43705\,
            I => \N__43649\
        );

    \I__10026\ : InMux
    port map (
            O => \N__43704\,
            I => \N__43649\
        );

    \I__10025\ : InMux
    port map (
            O => \N__43703\,
            I => \N__43649\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__43694\,
            I => \N__43634\
        );

    \I__10023\ : LocalMux
    port map (
            O => \N__43685\,
            I => \N__43634\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43634\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__43667\,
            I => \N__43634\
        );

    \I__10020\ : LocalMux
    port map (
            O => \N__43658\,
            I => \N__43629\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__43649\,
            I => \N__43629\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43648\,
            I => \N__43624\
        );

    \I__10017\ : InMux
    port map (
            O => \N__43647\,
            I => \N__43624\
        );

    \I__10016\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43615\
        );

    \I__10015\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43615\
        );

    \I__10014\ : InMux
    port map (
            O => \N__43644\,
            I => \N__43615\
        );

    \I__10013\ : InMux
    port map (
            O => \N__43643\,
            I => \N__43615\
        );

    \I__10012\ : Span4Mux_v
    port map (
            O => \N__43634\,
            I => \N__43606\
        );

    \I__10011\ : Span4Mux_v
    port map (
            O => \N__43629\,
            I => \N__43606\
        );

    \I__10010\ : LocalMux
    port map (
            O => \N__43624\,
            I => \N__43606\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43615\,
            I => \N__43606\
        );

    \I__10008\ : Span4Mux_h
    port map (
            O => \N__43606\,
            I => \N__43603\
        );

    \I__10007\ : Odrv4
    port map (
            O => \N__43603\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10006\ : InMux
    port map (
            O => \N__43600\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__10005\ : CascadeMux
    port map (
            O => \N__43597\,
            I => \N__43594\
        );

    \I__10004\ : InMux
    port map (
            O => \N__43594\,
            I => \N__43591\
        );

    \I__10003\ : LocalMux
    port map (
            O => \N__43591\,
            I => \N__43587\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43590\,
            I => \N__43584\
        );

    \I__10001\ : Span4Mux_v
    port map (
            O => \N__43587\,
            I => \N__43581\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__43584\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__9999\ : Odrv4
    port map (
            O => \N__43581\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__9998\ : CEMux
    port map (
            O => \N__43576\,
            I => \N__43573\
        );

    \I__9997\ : LocalMux
    port map (
            O => \N__43573\,
            I => \N__43568\
        );

    \I__9996\ : CEMux
    port map (
            O => \N__43572\,
            I => \N__43565\
        );

    \I__9995\ : CEMux
    port map (
            O => \N__43571\,
            I => \N__43562\
        );

    \I__9994\ : Span4Mux_v
    port map (
            O => \N__43568\,
            I => \N__43556\
        );

    \I__9993\ : LocalMux
    port map (
            O => \N__43565\,
            I => \N__43556\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__43562\,
            I => \N__43553\
        );

    \I__9991\ : CEMux
    port map (
            O => \N__43561\,
            I => \N__43550\
        );

    \I__9990\ : Span4Mux_v
    port map (
            O => \N__43556\,
            I => \N__43545\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__43553\,
            I => \N__43545\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__43550\,
            I => \N__43542\
        );

    \I__9987\ : Span4Mux_h
    port map (
            O => \N__43545\,
            I => \N__43539\
        );

    \I__9986\ : Span4Mux_h
    port map (
            O => \N__43542\,
            I => \N__43536\
        );

    \I__9985\ : Odrv4
    port map (
            O => \N__43539\,
            I => \current_shift_inst.timer_s1.N_191_i\
        );

    \I__9984\ : Odrv4
    port map (
            O => \N__43536\,
            I => \current_shift_inst.timer_s1.N_191_i\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43531\,
            I => \N__43528\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__43528\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\
        );

    \I__9981\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43522\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__43522\,
            I => \N__43519\
        );

    \I__9979\ : Odrv12
    port map (
            O => \N__43519\,
            I => \current_shift_inst.un4_control_input_axb_14\
        );

    \I__9978\ : InMux
    port map (
            O => \N__43516\,
            I => \N__43513\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__43513\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\
        );

    \I__9976\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43507\
        );

    \I__9975\ : LocalMux
    port map (
            O => \N__43507\,
            I => \N__43504\
        );

    \I__9974\ : Odrv12
    port map (
            O => \N__43504\,
            I => \current_shift_inst.un4_control_input_axb_24\
        );

    \I__9973\ : InMux
    port map (
            O => \N__43501\,
            I => \N__43490\
        );

    \I__9972\ : InMux
    port map (
            O => \N__43500\,
            I => \N__43483\
        );

    \I__9971\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43483\
        );

    \I__9970\ : InMux
    port map (
            O => \N__43498\,
            I => \N__43483\
        );

    \I__9969\ : InMux
    port map (
            O => \N__43497\,
            I => \N__43474\
        );

    \I__9968\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43474\
        );

    \I__9967\ : InMux
    port map (
            O => \N__43495\,
            I => \N__43474\
        );

    \I__9966\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43474\
        );

    \I__9965\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43446\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__43490\,
            I => \N__43443\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__43483\,
            I => \N__43438\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__43474\,
            I => \N__43438\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43473\,
            I => \N__43435\
        );

    \I__9960\ : CascadeMux
    port map (
            O => \N__43472\,
            I => \N__43431\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__43471\,
            I => \N__43427\
        );

    \I__9958\ : CascadeMux
    port map (
            O => \N__43470\,
            I => \N__43424\
        );

    \I__9957\ : CascadeMux
    port map (
            O => \N__43469\,
            I => \N__43421\
        );

    \I__9956\ : CascadeMux
    port map (
            O => \N__43468\,
            I => \N__43418\
        );

    \I__9955\ : CascadeMux
    port map (
            O => \N__43467\,
            I => \N__43415\
        );

    \I__9954\ : CascadeMux
    port map (
            O => \N__43466\,
            I => \N__43412\
        );

    \I__9953\ : CascadeMux
    port map (
            O => \N__43465\,
            I => \N__43409\
        );

    \I__9952\ : CascadeMux
    port map (
            O => \N__43464\,
            I => \N__43406\
        );

    \I__9951\ : CascadeMux
    port map (
            O => \N__43463\,
            I => \N__43403\
        );

    \I__9950\ : CascadeMux
    port map (
            O => \N__43462\,
            I => \N__43400\
        );

    \I__9949\ : CascadeMux
    port map (
            O => \N__43461\,
            I => \N__43397\
        );

    \I__9948\ : CascadeMux
    port map (
            O => \N__43460\,
            I => \N__43394\
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__43459\,
            I => \N__43391\
        );

    \I__9946\ : CascadeMux
    port map (
            O => \N__43458\,
            I => \N__43388\
        );

    \I__9945\ : CascadeMux
    port map (
            O => \N__43457\,
            I => \N__43385\
        );

    \I__9944\ : CascadeMux
    port map (
            O => \N__43456\,
            I => \N__43382\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__43455\,
            I => \N__43379\
        );

    \I__9942\ : CascadeMux
    port map (
            O => \N__43454\,
            I => \N__43376\
        );

    \I__9941\ : CascadeMux
    port map (
            O => \N__43453\,
            I => \N__43373\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__43452\,
            I => \N__43370\
        );

    \I__9939\ : CascadeMux
    port map (
            O => \N__43451\,
            I => \N__43367\
        );

    \I__9938\ : CascadeMux
    port map (
            O => \N__43450\,
            I => \N__43364\
        );

    \I__9937\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43354\
        );

    \I__9936\ : LocalMux
    port map (
            O => \N__43446\,
            I => \N__43351\
        );

    \I__9935\ : Span4Mux_h
    port map (
            O => \N__43443\,
            I => \N__43345\
        );

    \I__9934\ : Span4Mux_v
    port map (
            O => \N__43438\,
            I => \N__43345\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__43435\,
            I => \N__43342\
        );

    \I__9932\ : CascadeMux
    port map (
            O => \N__43434\,
            I => \N__43331\
        );

    \I__9931\ : InMux
    port map (
            O => \N__43431\,
            I => \N__43326\
        );

    \I__9930\ : InMux
    port map (
            O => \N__43430\,
            I => \N__43326\
        );

    \I__9929\ : InMux
    port map (
            O => \N__43427\,
            I => \N__43317\
        );

    \I__9928\ : InMux
    port map (
            O => \N__43424\,
            I => \N__43317\
        );

    \I__9927\ : InMux
    port map (
            O => \N__43421\,
            I => \N__43317\
        );

    \I__9926\ : InMux
    port map (
            O => \N__43418\,
            I => \N__43317\
        );

    \I__9925\ : InMux
    port map (
            O => \N__43415\,
            I => \N__43308\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43412\,
            I => \N__43308\
        );

    \I__9923\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43308\
        );

    \I__9922\ : InMux
    port map (
            O => \N__43406\,
            I => \N__43308\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43403\,
            I => \N__43301\
        );

    \I__9920\ : InMux
    port map (
            O => \N__43400\,
            I => \N__43301\
        );

    \I__9919\ : InMux
    port map (
            O => \N__43397\,
            I => \N__43301\
        );

    \I__9918\ : InMux
    port map (
            O => \N__43394\,
            I => \N__43294\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43294\
        );

    \I__9916\ : InMux
    port map (
            O => \N__43388\,
            I => \N__43294\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43385\,
            I => \N__43285\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43285\
        );

    \I__9913\ : InMux
    port map (
            O => \N__43379\,
            I => \N__43285\
        );

    \I__9912\ : InMux
    port map (
            O => \N__43376\,
            I => \N__43285\
        );

    \I__9911\ : InMux
    port map (
            O => \N__43373\,
            I => \N__43276\
        );

    \I__9910\ : InMux
    port map (
            O => \N__43370\,
            I => \N__43276\
        );

    \I__9909\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43276\
        );

    \I__9908\ : InMux
    port map (
            O => \N__43364\,
            I => \N__43276\
        );

    \I__9907\ : CascadeMux
    port map (
            O => \N__43363\,
            I => \N__43273\
        );

    \I__9906\ : CascadeMux
    port map (
            O => \N__43362\,
            I => \N__43270\
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__43361\,
            I => \N__43267\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__43360\,
            I => \N__43264\
        );

    \I__9903\ : CascadeMux
    port map (
            O => \N__43359\,
            I => \N__43261\
        );

    \I__9902\ : CascadeMux
    port map (
            O => \N__43358\,
            I => \N__43258\
        );

    \I__9901\ : CascadeMux
    port map (
            O => \N__43357\,
            I => \N__43255\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__43354\,
            I => \N__43250\
        );

    \I__9899\ : Span4Mux_s1_v
    port map (
            O => \N__43351\,
            I => \N__43250\
        );

    \I__9898\ : InMux
    port map (
            O => \N__43350\,
            I => \N__43247\
        );

    \I__9897\ : Span4Mux_v
    port map (
            O => \N__43345\,
            I => \N__43242\
        );

    \I__9896\ : Span4Mux_v
    port map (
            O => \N__43342\,
            I => \N__43242\
        );

    \I__9895\ : InMux
    port map (
            O => \N__43341\,
            I => \N__43235\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43340\,
            I => \N__43235\
        );

    \I__9893\ : InMux
    port map (
            O => \N__43339\,
            I => \N__43235\
        );

    \I__9892\ : InMux
    port map (
            O => \N__43338\,
            I => \N__43226\
        );

    \I__9891\ : InMux
    port map (
            O => \N__43337\,
            I => \N__43226\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43226\
        );

    \I__9889\ : InMux
    port map (
            O => \N__43335\,
            I => \N__43226\
        );

    \I__9888\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43223\
        );

    \I__9887\ : InMux
    port map (
            O => \N__43331\,
            I => \N__43220\
        );

    \I__9886\ : LocalMux
    port map (
            O => \N__43326\,
            I => \N__43217\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__43317\,
            I => \N__43212\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__43308\,
            I => \N__43212\
        );

    \I__9883\ : LocalMux
    port map (
            O => \N__43301\,
            I => \N__43203\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43294\,
            I => \N__43203\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43285\,
            I => \N__43203\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__43276\,
            I => \N__43203\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43196\
        );

    \I__9878\ : InMux
    port map (
            O => \N__43270\,
            I => \N__43196\
        );

    \I__9877\ : InMux
    port map (
            O => \N__43267\,
            I => \N__43196\
        );

    \I__9876\ : InMux
    port map (
            O => \N__43264\,
            I => \N__43187\
        );

    \I__9875\ : InMux
    port map (
            O => \N__43261\,
            I => \N__43187\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43258\,
            I => \N__43187\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43255\,
            I => \N__43187\
        );

    \I__9872\ : Sp12to4
    port map (
            O => \N__43250\,
            I => \N__43182\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43247\,
            I => \N__43182\
        );

    \I__9870\ : Span4Mux_h
    port map (
            O => \N__43242\,
            I => \N__43179\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__43235\,
            I => \N__43174\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__43226\,
            I => \N__43174\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__43223\,
            I => \N__43171\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__43220\,
            I => \N__43166\
        );

    \I__9865\ : Sp12to4
    port map (
            O => \N__43217\,
            I => \N__43166\
        );

    \I__9864\ : Span4Mux_v
    port map (
            O => \N__43212\,
            I => \N__43163\
        );

    \I__9863\ : Span4Mux_v
    port map (
            O => \N__43203\,
            I => \N__43156\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__43196\,
            I => \N__43156\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43187\,
            I => \N__43156\
        );

    \I__9860\ : Span12Mux_s7_h
    port map (
            O => \N__43182\,
            I => \N__43153\
        );

    \I__9859\ : Sp12to4
    port map (
            O => \N__43179\,
            I => \N__43148\
        );

    \I__9858\ : Span12Mux_s5_h
    port map (
            O => \N__43174\,
            I => \N__43148\
        );

    \I__9857\ : Span12Mux_s10_h
    port map (
            O => \N__43171\,
            I => \N__43145\
        );

    \I__9856\ : Span12Mux_v
    port map (
            O => \N__43166\,
            I => \N__43142\
        );

    \I__9855\ : Span4Mux_h
    port map (
            O => \N__43163\,
            I => \N__43137\
        );

    \I__9854\ : Span4Mux_h
    port map (
            O => \N__43156\,
            I => \N__43137\
        );

    \I__9853\ : Span12Mux_v
    port map (
            O => \N__43153\,
            I => \N__43134\
        );

    \I__9852\ : Span12Mux_h
    port map (
            O => \N__43148\,
            I => \N__43131\
        );

    \I__9851\ : Span12Mux_v
    port map (
            O => \N__43145\,
            I => \N__43126\
        );

    \I__9850\ : Span12Mux_h
    port map (
            O => \N__43142\,
            I => \N__43126\
        );

    \I__9849\ : Span4Mux_v
    port map (
            O => \N__43137\,
            I => \N__43123\
        );

    \I__9848\ : Odrv12
    port map (
            O => \N__43134\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9847\ : Odrv12
    port map (
            O => \N__43131\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9846\ : Odrv12
    port map (
            O => \N__43126\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9845\ : Odrv4
    port map (
            O => \N__43123\,
            I => \CONSTANT_ONE_NET\
        );

    \I__9844\ : CascadeMux
    port map (
            O => \N__43114\,
            I => \N__43110\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43113\,
            I => \N__43107\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43110\,
            I => \N__43104\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43107\,
            I => \N__43098\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__43104\,
            I => \N__43098\
        );

    \I__9839\ : InMux
    port map (
            O => \N__43103\,
            I => \N__43095\
        );

    \I__9838\ : Span4Mux_v
    port map (
            O => \N__43098\,
            I => \N__43092\
        );

    \I__9837\ : LocalMux
    port map (
            O => \N__43095\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9836\ : Odrv4
    port map (
            O => \N__43092\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43087\,
            I => \bfn_17_13_0_\
        );

    \I__9834\ : CascadeMux
    port map (
            O => \N__43084\,
            I => \N__43080\
        );

    \I__9833\ : InMux
    port map (
            O => \N__43083\,
            I => \N__43077\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43080\,
            I => \N__43074\
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__43077\,
            I => \N__43068\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__43074\,
            I => \N__43068\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43073\,
            I => \N__43065\
        );

    \I__9828\ : Span4Mux_v
    port map (
            O => \N__43068\,
            I => \N__43062\
        );

    \I__9827\ : LocalMux
    port map (
            O => \N__43065\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9826\ : Odrv4
    port map (
            O => \N__43062\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43057\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__9824\ : CascadeMux
    port map (
            O => \N__43054\,
            I => \N__43050\
        );

    \I__9823\ : CascadeMux
    port map (
            O => \N__43053\,
            I => \N__43047\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43050\,
            I => \N__43041\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43047\,
            I => \N__43041\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43046\,
            I => \N__43038\
        );

    \I__9819\ : LocalMux
    port map (
            O => \N__43041\,
            I => \N__43035\
        );

    \I__9818\ : LocalMux
    port map (
            O => \N__43038\,
            I => \N__43030\
        );

    \I__9817\ : Span4Mux_v
    port map (
            O => \N__43035\,
            I => \N__43030\
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__43030\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43027\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__9814\ : CascadeMux
    port map (
            O => \N__43024\,
            I => \N__43020\
        );

    \I__9813\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43016\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43020\,
            I => \N__43013\
        );

    \I__9811\ : InMux
    port map (
            O => \N__43019\,
            I => \N__43010\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43016\,
            I => \N__43005\
        );

    \I__9809\ : LocalMux
    port map (
            O => \N__43013\,
            I => \N__43005\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__43010\,
            I => \N__43000\
        );

    \I__9807\ : Span4Mux_v
    port map (
            O => \N__43005\,
            I => \N__43000\
        );

    \I__9806\ : Odrv4
    port map (
            O => \N__43000\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9805\ : InMux
    port map (
            O => \N__42997\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__9804\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42988\
        );

    \I__9803\ : InMux
    port map (
            O => \N__42993\,
            I => \N__42988\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__42988\,
            I => \N__42984\
        );

    \I__9801\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42981\
        );

    \I__9800\ : Span4Mux_v
    port map (
            O => \N__42984\,
            I => \N__42978\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__42981\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9798\ : Odrv4
    port map (
            O => \N__42978\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9797\ : InMux
    port map (
            O => \N__42973\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__9796\ : CascadeMux
    port map (
            O => \N__42970\,
            I => \N__42966\
        );

    \I__9795\ : CascadeMux
    port map (
            O => \N__42969\,
            I => \N__42963\
        );

    \I__9794\ : InMux
    port map (
            O => \N__42966\,
            I => \N__42958\
        );

    \I__9793\ : InMux
    port map (
            O => \N__42963\,
            I => \N__42958\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__42958\,
            I => \N__42954\
        );

    \I__9791\ : InMux
    port map (
            O => \N__42957\,
            I => \N__42951\
        );

    \I__9790\ : Span4Mux_v
    port map (
            O => \N__42954\,
            I => \N__42948\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__42951\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9788\ : Odrv4
    port map (
            O => \N__42948\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9787\ : InMux
    port map (
            O => \N__42943\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__9786\ : CascadeMux
    port map (
            O => \N__42940\,
            I => \N__42936\
        );

    \I__9785\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42933\
        );

    \I__9784\ : InMux
    port map (
            O => \N__42936\,
            I => \N__42930\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__42933\,
            I => \N__42924\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__42930\,
            I => \N__42924\
        );

    \I__9781\ : InMux
    port map (
            O => \N__42929\,
            I => \N__42921\
        );

    \I__9780\ : Span4Mux_v
    port map (
            O => \N__42924\,
            I => \N__42918\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__42921\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9778\ : Odrv4
    port map (
            O => \N__42918\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9777\ : InMux
    port map (
            O => \N__42913\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__9776\ : InMux
    port map (
            O => \N__42910\,
            I => \N__42904\
        );

    \I__9775\ : InMux
    port map (
            O => \N__42909\,
            I => \N__42904\
        );

    \I__9774\ : LocalMux
    port map (
            O => \N__42904\,
            I => \N__42900\
        );

    \I__9773\ : InMux
    port map (
            O => \N__42903\,
            I => \N__42897\
        );

    \I__9772\ : Span4Mux_v
    port map (
            O => \N__42900\,
            I => \N__42894\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__42897\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9770\ : Odrv4
    port map (
            O => \N__42894\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9769\ : InMux
    port map (
            O => \N__42889\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__9768\ : CascadeMux
    port map (
            O => \N__42886\,
            I => \N__42882\
        );

    \I__9767\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42879\
        );

    \I__9766\ : InMux
    port map (
            O => \N__42882\,
            I => \N__42876\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__42879\,
            I => \N__42870\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__42876\,
            I => \N__42870\
        );

    \I__9763\ : InMux
    port map (
            O => \N__42875\,
            I => \N__42867\
        );

    \I__9762\ : Span4Mux_v
    port map (
            O => \N__42870\,
            I => \N__42864\
        );

    \I__9761\ : LocalMux
    port map (
            O => \N__42867\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9760\ : Odrv4
    port map (
            O => \N__42864\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9759\ : CascadeMux
    port map (
            O => \N__42859\,
            I => \N__42855\
        );

    \I__9758\ : InMux
    port map (
            O => \N__42858\,
            I => \N__42852\
        );

    \I__9757\ : InMux
    port map (
            O => \N__42855\,
            I => \N__42849\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__42852\,
            I => \N__42843\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__42849\,
            I => \N__42843\
        );

    \I__9754\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42840\
        );

    \I__9753\ : Span4Mux_v
    port map (
            O => \N__42843\,
            I => \N__42837\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__42840\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9751\ : Odrv4
    port map (
            O => \N__42837\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9750\ : InMux
    port map (
            O => \N__42832\,
            I => \bfn_17_12_0_\
        );

    \I__9749\ : CascadeMux
    port map (
            O => \N__42829\,
            I => \N__42825\
        );

    \I__9748\ : CascadeMux
    port map (
            O => \N__42828\,
            I => \N__42822\
        );

    \I__9747\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42819\
        );

    \I__9746\ : InMux
    port map (
            O => \N__42822\,
            I => \N__42816\
        );

    \I__9745\ : LocalMux
    port map (
            O => \N__42819\,
            I => \N__42810\
        );

    \I__9744\ : LocalMux
    port map (
            O => \N__42816\,
            I => \N__42810\
        );

    \I__9743\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42807\
        );

    \I__9742\ : Span4Mux_v
    port map (
            O => \N__42810\,
            I => \N__42804\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__42807\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9740\ : Odrv4
    port map (
            O => \N__42804\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9739\ : InMux
    port map (
            O => \N__42799\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__9738\ : CascadeMux
    port map (
            O => \N__42796\,
            I => \N__42792\
        );

    \I__9737\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42788\
        );

    \I__9736\ : InMux
    port map (
            O => \N__42792\,
            I => \N__42785\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42791\,
            I => \N__42782\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__42788\,
            I => \N__42777\
        );

    \I__9733\ : LocalMux
    port map (
            O => \N__42785\,
            I => \N__42777\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__42782\,
            I => \N__42772\
        );

    \I__9731\ : Span4Mux_v
    port map (
            O => \N__42777\,
            I => \N__42772\
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__42772\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__9729\ : InMux
    port map (
            O => \N__42769\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__9728\ : InMux
    port map (
            O => \N__42766\,
            I => \N__42759\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42759\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42764\,
            I => \N__42756\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__42759\,
            I => \N__42753\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__42756\,
            I => \N__42748\
        );

    \I__9723\ : Span4Mux_v
    port map (
            O => \N__42753\,
            I => \N__42748\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__42748\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__9721\ : InMux
    port map (
            O => \N__42745\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__42742\,
            I => \N__42738\
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__42741\,
            I => \N__42735\
        );

    \I__9718\ : InMux
    port map (
            O => \N__42738\,
            I => \N__42730\
        );

    \I__9717\ : InMux
    port map (
            O => \N__42735\,
            I => \N__42730\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__42730\,
            I => \N__42726\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42729\,
            I => \N__42723\
        );

    \I__9714\ : Span4Mux_v
    port map (
            O => \N__42726\,
            I => \N__42720\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__42723\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__9712\ : Odrv4
    port map (
            O => \N__42720\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__9711\ : InMux
    port map (
            O => \N__42715\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__9710\ : CascadeMux
    port map (
            O => \N__42712\,
            I => \N__42708\
        );

    \I__9709\ : CascadeMux
    port map (
            O => \N__42711\,
            I => \N__42705\
        );

    \I__9708\ : InMux
    port map (
            O => \N__42708\,
            I => \N__42700\
        );

    \I__9707\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42700\
        );

    \I__9706\ : LocalMux
    port map (
            O => \N__42700\,
            I => \N__42696\
        );

    \I__9705\ : InMux
    port map (
            O => \N__42699\,
            I => \N__42693\
        );

    \I__9704\ : Span4Mux_v
    port map (
            O => \N__42696\,
            I => \N__42690\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__42693\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__9702\ : Odrv4
    port map (
            O => \N__42690\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42685\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42682\,
            I => \N__42676\
        );

    \I__9699\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42676\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__42676\,
            I => \N__42672\
        );

    \I__9697\ : InMux
    port map (
            O => \N__42675\,
            I => \N__42669\
        );

    \I__9696\ : Span4Mux_v
    port map (
            O => \N__42672\,
            I => \N__42666\
        );

    \I__9695\ : LocalMux
    port map (
            O => \N__42669\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__9694\ : Odrv4
    port map (
            O => \N__42666\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__9693\ : InMux
    port map (
            O => \N__42661\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__9692\ : InMux
    port map (
            O => \N__42658\,
            I => \N__42652\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42657\,
            I => \N__42652\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__42652\,
            I => \N__42648\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42651\,
            I => \N__42645\
        );

    \I__9688\ : Span4Mux_v
    port map (
            O => \N__42648\,
            I => \N__42642\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__42645\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9686\ : Odrv4
    port map (
            O => \N__42642\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42637\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__9684\ : CascadeMux
    port map (
            O => \N__42634\,
            I => \N__42631\
        );

    \I__9683\ : InMux
    port map (
            O => \N__42631\,
            I => \N__42623\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42630\,
            I => \N__42623\
        );

    \I__9681\ : InMux
    port map (
            O => \N__42629\,
            I => \N__42618\
        );

    \I__9680\ : InMux
    port map (
            O => \N__42628\,
            I => \N__42618\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__42623\,
            I => \N__42615\
        );

    \I__9678\ : LocalMux
    port map (
            O => \N__42618\,
            I => \N__42612\
        );

    \I__9677\ : Span4Mux_v
    port map (
            O => \N__42615\,
            I => \N__42609\
        );

    \I__9676\ : Span4Mux_v
    port map (
            O => \N__42612\,
            I => \N__42606\
        );

    \I__9675\ : Odrv4
    port map (
            O => \N__42609\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__42606\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__9673\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42595\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42600\,
            I => \N__42595\
        );

    \I__9671\ : LocalMux
    port map (
            O => \N__42595\,
            I => \N__42592\
        );

    \I__9670\ : Span4Mux_v
    port map (
            O => \N__42592\,
            I => \N__42585\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42591\,
            I => \N__42580\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42590\,
            I => \N__42580\
        );

    \I__9667\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42575\
        );

    \I__9666\ : InMux
    port map (
            O => \N__42588\,
            I => \N__42575\
        );

    \I__9665\ : Odrv4
    port map (
            O => \N__42585\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__42580\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__42575\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__9662\ : InMux
    port map (
            O => \N__42568\,
            I => \N__42564\
        );

    \I__9661\ : CascadeMux
    port map (
            O => \N__42567\,
            I => \N__42561\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__42564\,
            I => \N__42558\
        );

    \I__9659\ : InMux
    port map (
            O => \N__42561\,
            I => \N__42555\
        );

    \I__9658\ : Span4Mux_h
    port map (
            O => \N__42558\,
            I => \N__42549\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__42555\,
            I => \N__42549\
        );

    \I__9656\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42546\
        );

    \I__9655\ : Span4Mux_v
    port map (
            O => \N__42549\,
            I => \N__42543\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__42546\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9653\ : Odrv4
    port map (
            O => \N__42543\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9652\ : InMux
    port map (
            O => \N__42538\,
            I => \bfn_17_11_0_\
        );

    \I__9651\ : InMux
    port map (
            O => \N__42535\,
            I => \N__42532\
        );

    \I__9650\ : LocalMux
    port map (
            O => \N__42532\,
            I => \N__42528\
        );

    \I__9649\ : CascadeMux
    port map (
            O => \N__42531\,
            I => \N__42525\
        );

    \I__9648\ : Span4Mux_h
    port map (
            O => \N__42528\,
            I => \N__42522\
        );

    \I__9647\ : InMux
    port map (
            O => \N__42525\,
            I => \N__42519\
        );

    \I__9646\ : Span4Mux_h
    port map (
            O => \N__42522\,
            I => \N__42513\
        );

    \I__9645\ : LocalMux
    port map (
            O => \N__42519\,
            I => \N__42513\
        );

    \I__9644\ : InMux
    port map (
            O => \N__42518\,
            I => \N__42510\
        );

    \I__9643\ : Span4Mux_v
    port map (
            O => \N__42513\,
            I => \N__42507\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__42510\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9641\ : Odrv4
    port map (
            O => \N__42507\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9640\ : InMux
    port map (
            O => \N__42502\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42499\,
            I => \N__42492\
        );

    \I__9638\ : InMux
    port map (
            O => \N__42498\,
            I => \N__42492\
        );

    \I__9637\ : InMux
    port map (
            O => \N__42497\,
            I => \N__42489\
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__42492\,
            I => \N__42486\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__42489\,
            I => \N__42481\
        );

    \I__9634\ : Span4Mux_v
    port map (
            O => \N__42486\,
            I => \N__42481\
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__42481\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9632\ : InMux
    port map (
            O => \N__42478\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__9631\ : InMux
    port map (
            O => \N__42475\,
            I => \N__42469\
        );

    \I__9630\ : InMux
    port map (
            O => \N__42474\,
            I => \N__42469\
        );

    \I__9629\ : LocalMux
    port map (
            O => \N__42469\,
            I => \N__42465\
        );

    \I__9628\ : InMux
    port map (
            O => \N__42468\,
            I => \N__42462\
        );

    \I__9627\ : Sp12to4
    port map (
            O => \N__42465\,
            I => \N__42459\
        );

    \I__9626\ : LocalMux
    port map (
            O => \N__42462\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9625\ : Odrv12
    port map (
            O => \N__42459\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9624\ : InMux
    port map (
            O => \N__42454\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__9623\ : CascadeMux
    port map (
            O => \N__42451\,
            I => \N__42447\
        );

    \I__9622\ : CascadeMux
    port map (
            O => \N__42450\,
            I => \N__42444\
        );

    \I__9621\ : InMux
    port map (
            O => \N__42447\,
            I => \N__42439\
        );

    \I__9620\ : InMux
    port map (
            O => \N__42444\,
            I => \N__42439\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__42439\,
            I => \N__42435\
        );

    \I__9618\ : InMux
    port map (
            O => \N__42438\,
            I => \N__42432\
        );

    \I__9617\ : Span4Mux_v
    port map (
            O => \N__42435\,
            I => \N__42429\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__42432\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9615\ : Odrv4
    port map (
            O => \N__42429\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9614\ : InMux
    port map (
            O => \N__42424\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__9613\ : CascadeMux
    port map (
            O => \N__42421\,
            I => \N__42417\
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__42420\,
            I => \N__42414\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42417\,
            I => \N__42409\
        );

    \I__9610\ : InMux
    port map (
            O => \N__42414\,
            I => \N__42409\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__42409\,
            I => \N__42405\
        );

    \I__9608\ : InMux
    port map (
            O => \N__42408\,
            I => \N__42402\
        );

    \I__9607\ : Span4Mux_v
    port map (
            O => \N__42405\,
            I => \N__42399\
        );

    \I__9606\ : LocalMux
    port map (
            O => \N__42402\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9605\ : Odrv4
    port map (
            O => \N__42399\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42394\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__9603\ : InMux
    port map (
            O => \N__42391\,
            I => \N__42385\
        );

    \I__9602\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42385\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__42385\,
            I => \N__42381\
        );

    \I__9600\ : InMux
    port map (
            O => \N__42384\,
            I => \N__42378\
        );

    \I__9599\ : Span4Mux_v
    port map (
            O => \N__42381\,
            I => \N__42375\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__42378\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9597\ : Odrv4
    port map (
            O => \N__42375\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42370\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42367\,
            I => \N__42361\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42366\,
            I => \N__42361\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__42361\,
            I => \N__42357\
        );

    \I__9592\ : InMux
    port map (
            O => \N__42360\,
            I => \N__42354\
        );

    \I__9591\ : Span4Mux_v
    port map (
            O => \N__42357\,
            I => \N__42351\
        );

    \I__9590\ : LocalMux
    port map (
            O => \N__42354\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9589\ : Odrv4
    port map (
            O => \N__42351\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9588\ : InMux
    port map (
            O => \N__42346\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__9587\ : InMux
    port map (
            O => \N__42343\,
            I => \N__42340\
        );

    \I__9586\ : LocalMux
    port map (
            O => \N__42340\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__9585\ : CascadeMux
    port map (
            O => \N__42337\,
            I => \phase_controller_slave.N_214_cascade_\
        );

    \I__9584\ : CascadeMux
    port map (
            O => \N__42334\,
            I => \N__42328\
        );

    \I__9583\ : CascadeMux
    port map (
            O => \N__42333\,
            I => \N__42325\
        );

    \I__9582\ : CascadeMux
    port map (
            O => \N__42332\,
            I => \N__42322\
        );

    \I__9581\ : CascadeMux
    port map (
            O => \N__42331\,
            I => \N__42319\
        );

    \I__9580\ : InMux
    port map (
            O => \N__42328\,
            I => \N__42296\
        );

    \I__9579\ : InMux
    port map (
            O => \N__42325\,
            I => \N__42296\
        );

    \I__9578\ : InMux
    port map (
            O => \N__42322\,
            I => \N__42296\
        );

    \I__9577\ : InMux
    port map (
            O => \N__42319\,
            I => \N__42296\
        );

    \I__9576\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42287\
        );

    \I__9575\ : InMux
    port map (
            O => \N__42317\,
            I => \N__42287\
        );

    \I__9574\ : InMux
    port map (
            O => \N__42316\,
            I => \N__42287\
        );

    \I__9573\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42287\
        );

    \I__9572\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42272\
        );

    \I__9571\ : InMux
    port map (
            O => \N__42313\,
            I => \N__42272\
        );

    \I__9570\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42272\
        );

    \I__9569\ : InMux
    port map (
            O => \N__42311\,
            I => \N__42272\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42272\
        );

    \I__9567\ : InMux
    port map (
            O => \N__42309\,
            I => \N__42272\
        );

    \I__9566\ : InMux
    port map (
            O => \N__42308\,
            I => \N__42272\
        );

    \I__9565\ : CascadeMux
    port map (
            O => \N__42307\,
            I => \N__42267\
        );

    \I__9564\ : CascadeMux
    port map (
            O => \N__42306\,
            I => \N__42264\
        );

    \I__9563\ : InMux
    port map (
            O => \N__42305\,
            I => \N__42261\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__42296\,
            I => \N__42254\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__42287\,
            I => \N__42254\
        );

    \I__9560\ : LocalMux
    port map (
            O => \N__42272\,
            I => \N__42254\
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__42271\,
            I => \N__42251\
        );

    \I__9558\ : InMux
    port map (
            O => \N__42270\,
            I => \N__42247\
        );

    \I__9557\ : InMux
    port map (
            O => \N__42267\,
            I => \N__42242\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42264\,
            I => \N__42242\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__42261\,
            I => \N__42237\
        );

    \I__9554\ : Span4Mux_v
    port map (
            O => \N__42254\,
            I => \N__42237\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42251\,
            I => \N__42232\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42250\,
            I => \N__42232\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__42247\,
            I => \N__42227\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__42242\,
            I => \N__42220\
        );

    \I__9549\ : Span4Mux_h
    port map (
            O => \N__42237\,
            I => \N__42220\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__42232\,
            I => \N__42220\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42214\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42214\
        );

    \I__9545\ : Span4Mux_v
    port map (
            O => \N__42227\,
            I => \N__42211\
        );

    \I__9544\ : Span4Mux_h
    port map (
            O => \N__42220\,
            I => \N__42208\
        );

    \I__9543\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42205\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__42214\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9541\ : Odrv4
    port map (
            O => \N__42211\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9540\ : Odrv4
    port map (
            O => \N__42208\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__42205\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__9538\ : CascadeMux
    port map (
            O => \N__42196\,
            I => \N__42192\
        );

    \I__9537\ : CascadeMux
    port map (
            O => \N__42195\,
            I => \N__42184\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42179\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42179\
        );

    \I__9534\ : CascadeMux
    port map (
            O => \N__42190\,
            I => \N__42169\
        );

    \I__9533\ : CascadeMux
    port map (
            O => \N__42189\,
            I => \N__42166\
        );

    \I__9532\ : CascadeMux
    port map (
            O => \N__42188\,
            I => \N__42163\
        );

    \I__9531\ : CascadeMux
    port map (
            O => \N__42187\,
            I => \N__42160\
        );

    \I__9530\ : InMux
    port map (
            O => \N__42184\,
            I => \N__42157\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__42179\,
            I => \N__42154\
        );

    \I__9528\ : CascadeMux
    port map (
            O => \N__42178\,
            I => \N__42147\
        );

    \I__9527\ : CascadeMux
    port map (
            O => \N__42177\,
            I => \N__42144\
        );

    \I__9526\ : CascadeMux
    port map (
            O => \N__42176\,
            I => \N__42141\
        );

    \I__9525\ : CascadeMux
    port map (
            O => \N__42175\,
            I => \N__42138\
        );

    \I__9524\ : InMux
    port map (
            O => \N__42174\,
            I => \N__42117\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42173\,
            I => \N__42117\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42172\,
            I => \N__42117\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42117\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42166\,
            I => \N__42117\
        );

    \I__9519\ : InMux
    port map (
            O => \N__42163\,
            I => \N__42117\
        );

    \I__9518\ : InMux
    port map (
            O => \N__42160\,
            I => \N__42117\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42157\,
            I => \N__42114\
        );

    \I__9516\ : Span4Mux_h
    port map (
            O => \N__42154\,
            I => \N__42111\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42153\,
            I => \N__42102\
        );

    \I__9514\ : InMux
    port map (
            O => \N__42152\,
            I => \N__42102\
        );

    \I__9513\ : InMux
    port map (
            O => \N__42151\,
            I => \N__42102\
        );

    \I__9512\ : InMux
    port map (
            O => \N__42150\,
            I => \N__42102\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42147\,
            I => \N__42085\
        );

    \I__9510\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42085\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42141\,
            I => \N__42085\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42138\,
            I => \N__42085\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42085\
        );

    \I__9506\ : InMux
    port map (
            O => \N__42136\,
            I => \N__42085\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42085\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42134\,
            I => \N__42085\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42133\,
            I => \N__42080\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42132\,
            I => \N__42080\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42117\,
            I => \N__42077\
        );

    \I__9500\ : Span4Mux_v
    port map (
            O => \N__42114\,
            I => \N__42070\
        );

    \I__9499\ : Span4Mux_v
    port map (
            O => \N__42111\,
            I => \N__42070\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__42070\
        );

    \I__9497\ : LocalMux
    port map (
            O => \N__42085\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42080\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9495\ : Odrv4
    port map (
            O => \N__42077\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9494\ : Odrv4
    port map (
            O => \N__42070\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__9493\ : CascadeMux
    port map (
            O => \N__42061\,
            I => \N__42058\
        );

    \I__9492\ : InMux
    port map (
            O => \N__42058\,
            I => \N__42039\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42057\,
            I => \N__42024\
        );

    \I__9490\ : InMux
    port map (
            O => \N__42056\,
            I => \N__42024\
        );

    \I__9489\ : InMux
    port map (
            O => \N__42055\,
            I => \N__42024\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42024\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42024\
        );

    \I__9486\ : InMux
    port map (
            O => \N__42052\,
            I => \N__42024\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42051\,
            I => \N__42024\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42050\,
            I => \N__42007\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42049\,
            I => \N__42007\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42048\,
            I => \N__42007\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42047\,
            I => \N__42007\
        );

    \I__9480\ : InMux
    port map (
            O => \N__42046\,
            I => \N__42007\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42007\
        );

    \I__9478\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42007\
        );

    \I__9477\ : InMux
    port map (
            O => \N__42043\,
            I => \N__42007\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42042\,
            I => \N__41999\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42039\,
            I => \N__41994\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__42024\,
            I => \N__41994\
        );

    \I__9473\ : LocalMux
    port map (
            O => \N__42007\,
            I => \N__41991\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42006\,
            I => \N__41982\
        );

    \I__9471\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41982\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41982\
        );

    \I__9469\ : InMux
    port map (
            O => \N__42003\,
            I => \N__41982\
        );

    \I__9468\ : CascadeMux
    port map (
            O => \N__42002\,
            I => \N__41979\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__41999\,
            I => \N__41975\
        );

    \I__9466\ : Span4Mux_v
    port map (
            O => \N__41994\,
            I => \N__41968\
        );

    \I__9465\ : Span4Mux_v
    port map (
            O => \N__41991\,
            I => \N__41968\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__41982\,
            I => \N__41968\
        );

    \I__9463\ : InMux
    port map (
            O => \N__41979\,
            I => \N__41962\
        );

    \I__9462\ : InMux
    port map (
            O => \N__41978\,
            I => \N__41962\
        );

    \I__9461\ : Span4Mux_v
    port map (
            O => \N__41975\,
            I => \N__41959\
        );

    \I__9460\ : Span4Mux_h
    port map (
            O => \N__41968\,
            I => \N__41956\
        );

    \I__9459\ : InMux
    port map (
            O => \N__41967\,
            I => \N__41953\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__41962\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__41959\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__9456\ : Odrv4
    port map (
            O => \N__41956\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__41953\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__9454\ : CascadeMux
    port map (
            O => \N__41944\,
            I => \N__41941\
        );

    \I__9453\ : InMux
    port map (
            O => \N__41941\,
            I => \N__41938\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__41938\,
            I => \N__41935\
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__41935\,
            I => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__9450\ : CascadeMux
    port map (
            O => \N__41932\,
            I => \N__41928\
        );

    \I__9449\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41924\
        );

    \I__9448\ : InMux
    port map (
            O => \N__41928\,
            I => \N__41921\
        );

    \I__9447\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41918\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__41924\,
            I => \N__41913\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__41921\,
            I => \N__41913\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__41918\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__9443\ : Odrv4
    port map (
            O => \N__41913\,
            I => \current_shift_inst.timer_phase.counterZ0Z_27\
        );

    \I__9442\ : CascadeMux
    port map (
            O => \N__41908\,
            I => \N__41905\
        );

    \I__9441\ : InMux
    port map (
            O => \N__41905\,
            I => \N__41901\
        );

    \I__9440\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41898\
        );

    \I__9439\ : LocalMux
    port map (
            O => \N__41901\,
            I => \N__41895\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__41898\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__9437\ : Odrv4
    port map (
            O => \N__41895\,
            I => \current_shift_inst.timer_phase.counterZ0Z_29\
        );

    \I__9436\ : InMux
    port map (
            O => \N__41890\,
            I => \N__41887\
        );

    \I__9435\ : LocalMux
    port map (
            O => \N__41887\,
            I => \N__41883\
        );

    \I__9434\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41880\
        );

    \I__9433\ : Span4Mux_h
    port map (
            O => \N__41883\,
            I => \N__41877\
        );

    \I__9432\ : LocalMux
    port map (
            O => \N__41880\,
            I => \N__41874\
        );

    \I__9431\ : Span4Mux_v
    port map (
            O => \N__41877\,
            I => \N__41870\
        );

    \I__9430\ : Span12Mux_h
    port map (
            O => \N__41874\,
            I => \N__41867\
        );

    \I__9429\ : InMux
    port map (
            O => \N__41873\,
            I => \N__41864\
        );

    \I__9428\ : Odrv4
    port map (
            O => \N__41870\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__9427\ : Odrv12
    port map (
            O => \N__41867\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__41864\,
            I => \current_shift_inst.elapsed_time_ns_phase_30\
        );

    \I__9425\ : InMux
    port map (
            O => \N__41857\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\
        );

    \I__9424\ : InMux
    port map (
            O => \N__41854\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\
        );

    \I__9423\ : CascadeMux
    port map (
            O => \N__41851\,
            I => \N__41848\
        );

    \I__9422\ : InMux
    port map (
            O => \N__41848\,
            I => \N__41844\
        );

    \I__9421\ : CascadeMux
    port map (
            O => \N__41847\,
            I => \N__41841\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__41844\,
            I => \N__41838\
        );

    \I__9419\ : InMux
    port map (
            O => \N__41841\,
            I => \N__41835\
        );

    \I__9418\ : Span4Mux_h
    port map (
            O => \N__41838\,
            I => \N__41832\
        );

    \I__9417\ : LocalMux
    port map (
            O => \N__41835\,
            I => \N__41829\
        );

    \I__9416\ : Span4Mux_v
    port map (
            O => \N__41832\,
            I => \N__41824\
        );

    \I__9415\ : Span4Mux_h
    port map (
            O => \N__41829\,
            I => \N__41824\
        );

    \I__9414\ : Odrv4
    port map (
            O => \N__41824\,
            I => \current_shift_inst.elapsed_time_ns_phase_31\
        );

    \I__9413\ : CEMux
    port map (
            O => \N__41821\,
            I => \N__41806\
        );

    \I__9412\ : CEMux
    port map (
            O => \N__41820\,
            I => \N__41806\
        );

    \I__9411\ : CEMux
    port map (
            O => \N__41819\,
            I => \N__41806\
        );

    \I__9410\ : CEMux
    port map (
            O => \N__41818\,
            I => \N__41806\
        );

    \I__9409\ : CEMux
    port map (
            O => \N__41817\,
            I => \N__41806\
        );

    \I__9408\ : GlobalMux
    port map (
            O => \N__41806\,
            I => \N__41803\
        );

    \I__9407\ : gio2CtrlBuf
    port map (
            O => \N__41803\,
            I => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \I__9406\ : CascadeMux
    port map (
            O => \N__41800\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_\
        );

    \I__9405\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41794\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__41794\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\
        );

    \I__9403\ : InMux
    port map (
            O => \N__41791\,
            I => \N__41788\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__41788\,
            I => \N__41785\
        );

    \I__9401\ : Odrv4
    port map (
            O => \N__41785\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19\
        );

    \I__9400\ : InMux
    port map (
            O => \N__41782\,
            I => \N__41779\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__41779\,
            I => \N__41776\
        );

    \I__9398\ : Span4Mux_h
    port map (
            O => \N__41776\,
            I => \N__41773\
        );

    \I__9397\ : Span4Mux_h
    port map (
            O => \N__41773\,
            I => \N__41770\
        );

    \I__9396\ : Odrv4
    port map (
            O => \N__41770\,
            I => \il_max_comp2_D1\
        );

    \I__9395\ : InMux
    port map (
            O => \N__41767\,
            I => \N__41764\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__41764\,
            I => \N__41761\
        );

    \I__9393\ : Span4Mux_h
    port map (
            O => \N__41761\,
            I => \N__41758\
        );

    \I__9392\ : Span4Mux_h
    port map (
            O => \N__41758\,
            I => \N__41755\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__41755\,
            I => \il_min_comp2_D1\
        );

    \I__9390\ : CascadeMux
    port map (
            O => \N__41752\,
            I => \N__41747\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41744\
        );

    \I__9388\ : InMux
    port map (
            O => \N__41750\,
            I => \N__41741\
        );

    \I__9387\ : InMux
    port map (
            O => \N__41747\,
            I => \N__41738\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__41744\,
            I => \N__41731\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__41741\,
            I => \N__41731\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__41738\,
            I => \N__41731\
        );

    \I__9383\ : Odrv4
    port map (
            O => \N__41731\,
            I => \current_shift_inst.timer_phase.counterZ0Z_19\
        );

    \I__9382\ : InMux
    port map (
            O => \N__41728\,
            I => \N__41722\
        );

    \I__9381\ : InMux
    port map (
            O => \N__41727\,
            I => \N__41722\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__41722\,
            I => \N__41718\
        );

    \I__9379\ : InMux
    port map (
            O => \N__41721\,
            I => \N__41715\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__41718\,
            I => \N__41712\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__41715\,
            I => \N__41709\
        );

    \I__9376\ : Span4Mux_v
    port map (
            O => \N__41712\,
            I => \N__41706\
        );

    \I__9375\ : Span12Mux_v
    port map (
            O => \N__41709\,
            I => \N__41702\
        );

    \I__9374\ : Span4Mux_h
    port map (
            O => \N__41706\,
            I => \N__41699\
        );

    \I__9373\ : InMux
    port map (
            O => \N__41705\,
            I => \N__41696\
        );

    \I__9372\ : Odrv12
    port map (
            O => \N__41702\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__9371\ : Odrv4
    port map (
            O => \N__41699\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__41696\,
            I => \current_shift_inst.elapsed_time_ns_phase_22\
        );

    \I__9369\ : InMux
    port map (
            O => \N__41689\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\
        );

    \I__9368\ : CascadeMux
    port map (
            O => \N__41686\,
            I => \N__41682\
        );

    \I__9367\ : CascadeMux
    port map (
            O => \N__41685\,
            I => \N__41679\
        );

    \I__9366\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41673\
        );

    \I__9365\ : InMux
    port map (
            O => \N__41679\,
            I => \N__41673\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41678\,
            I => \N__41670\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__41673\,
            I => \N__41667\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41670\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__9361\ : Odrv4
    port map (
            O => \N__41667\,
            I => \current_shift_inst.timer_phase.counterZ0Z_20\
        );

    \I__9360\ : InMux
    port map (
            O => \N__41662\,
            I => \N__41658\
        );

    \I__9359\ : CascadeMux
    port map (
            O => \N__41661\,
            I => \N__41655\
        );

    \I__9358\ : LocalMux
    port map (
            O => \N__41658\,
            I => \N__41651\
        );

    \I__9357\ : InMux
    port map (
            O => \N__41655\,
            I => \N__41648\
        );

    \I__9356\ : InMux
    port map (
            O => \N__41654\,
            I => \N__41645\
        );

    \I__9355\ : Span4Mux_h
    port map (
            O => \N__41651\,
            I => \N__41642\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__41648\,
            I => \N__41639\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41645\,
            I => \N__41635\
        );

    \I__9352\ : Span4Mux_v
    port map (
            O => \N__41642\,
            I => \N__41632\
        );

    \I__9351\ : Span12Mux_h
    port map (
            O => \N__41639\,
            I => \N__41629\
        );

    \I__9350\ : InMux
    port map (
            O => \N__41638\,
            I => \N__41626\
        );

    \I__9349\ : Odrv12
    port map (
            O => \N__41635\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__9348\ : Odrv4
    port map (
            O => \N__41632\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__9347\ : Odrv12
    port map (
            O => \N__41629\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__41626\,
            I => \current_shift_inst.elapsed_time_ns_phase_23\
        );

    \I__9345\ : InMux
    port map (
            O => \N__41617\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\
        );

    \I__9344\ : CascadeMux
    port map (
            O => \N__41614\,
            I => \N__41610\
        );

    \I__9343\ : CascadeMux
    port map (
            O => \N__41613\,
            I => \N__41607\
        );

    \I__9342\ : InMux
    port map (
            O => \N__41610\,
            I => \N__41601\
        );

    \I__9341\ : InMux
    port map (
            O => \N__41607\,
            I => \N__41601\
        );

    \I__9340\ : InMux
    port map (
            O => \N__41606\,
            I => \N__41598\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__41601\,
            I => \N__41595\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__41598\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__9337\ : Odrv4
    port map (
            O => \N__41595\,
            I => \current_shift_inst.timer_phase.counterZ0Z_21\
        );

    \I__9336\ : CascadeMux
    port map (
            O => \N__41590\,
            I => \N__41587\
        );

    \I__9335\ : InMux
    port map (
            O => \N__41587\,
            I => \N__41584\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__41584\,
            I => \N__41581\
        );

    \I__9333\ : Span4Mux_h
    port map (
            O => \N__41581\,
            I => \N__41576\
        );

    \I__9332\ : InMux
    port map (
            O => \N__41580\,
            I => \N__41571\
        );

    \I__9331\ : InMux
    port map (
            O => \N__41579\,
            I => \N__41571\
        );

    \I__9330\ : Span4Mux_v
    port map (
            O => \N__41576\,
            I => \N__41567\
        );

    \I__9329\ : LocalMux
    port map (
            O => \N__41571\,
            I => \N__41564\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41570\,
            I => \N__41561\
        );

    \I__9327\ : Odrv4
    port map (
            O => \N__41567\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__9326\ : Odrv12
    port map (
            O => \N__41564\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__41561\,
            I => \current_shift_inst.elapsed_time_ns_phase_24\
        );

    \I__9324\ : InMux
    port map (
            O => \N__41554\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__41551\,
            I => \N__41548\
        );

    \I__9322\ : InMux
    port map (
            O => \N__41548\,
            I => \N__41543\
        );

    \I__9321\ : InMux
    port map (
            O => \N__41547\,
            I => \N__41540\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41546\,
            I => \N__41537\
        );

    \I__9319\ : LocalMux
    port map (
            O => \N__41543\,
            I => \N__41532\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__41540\,
            I => \N__41532\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41537\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__9316\ : Odrv12
    port map (
            O => \N__41532\,
            I => \current_shift_inst.timer_phase.counterZ0Z_22\
        );

    \I__9315\ : InMux
    port map (
            O => \N__41527\,
            I => \N__41521\
        );

    \I__9314\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41521\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__41521\,
            I => \N__41517\
        );

    \I__9312\ : InMux
    port map (
            O => \N__41520\,
            I => \N__41514\
        );

    \I__9311\ : Span4Mux_h
    port map (
            O => \N__41517\,
            I => \N__41511\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__41514\,
            I => \N__41507\
        );

    \I__9309\ : Span4Mux_v
    port map (
            O => \N__41511\,
            I => \N__41504\
        );

    \I__9308\ : InMux
    port map (
            O => \N__41510\,
            I => \N__41501\
        );

    \I__9307\ : Odrv12
    port map (
            O => \N__41507\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__9306\ : Odrv4
    port map (
            O => \N__41504\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__9305\ : LocalMux
    port map (
            O => \N__41501\,
            I => \current_shift_inst.elapsed_time_ns_phase_25\
        );

    \I__9304\ : InMux
    port map (
            O => \N__41494\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\
        );

    \I__9303\ : InMux
    port map (
            O => \N__41491\,
            I => \N__41485\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41490\,
            I => \N__41485\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__41485\,
            I => \N__41481\
        );

    \I__9300\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41478\
        );

    \I__9299\ : Span4Mux_h
    port map (
            O => \N__41481\,
            I => \N__41475\
        );

    \I__9298\ : LocalMux
    port map (
            O => \N__41478\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__41475\,
            I => \current_shift_inst.timer_phase.counterZ0Z_23\
        );

    \I__9296\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41465\
        );

    \I__9295\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41460\
        );

    \I__9294\ : InMux
    port map (
            O => \N__41468\,
            I => \N__41460\
        );

    \I__9293\ : LocalMux
    port map (
            O => \N__41465\,
            I => \N__41457\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__41460\,
            I => \N__41454\
        );

    \I__9291\ : Span4Mux_h
    port map (
            O => \N__41457\,
            I => \N__41451\
        );

    \I__9290\ : Span12Mux_v
    port map (
            O => \N__41454\,
            I => \N__41447\
        );

    \I__9289\ : Span4Mux_v
    port map (
            O => \N__41451\,
            I => \N__41444\
        );

    \I__9288\ : InMux
    port map (
            O => \N__41450\,
            I => \N__41441\
        );

    \I__9287\ : Odrv12
    port map (
            O => \N__41447\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__9286\ : Odrv4
    port map (
            O => \N__41444\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__41441\,
            I => \current_shift_inst.elapsed_time_ns_phase_26\
        );

    \I__9284\ : InMux
    port map (
            O => \N__41434\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\
        );

    \I__9283\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41427\
        );

    \I__9282\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41423\
        );

    \I__9281\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41420\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41426\,
            I => \N__41417\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__41423\,
            I => \N__41412\
        );

    \I__9278\ : Span4Mux_v
    port map (
            O => \N__41420\,
            I => \N__41412\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__41417\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__9276\ : Odrv4
    port map (
            O => \N__41412\,
            I => \current_shift_inst.timer_phase.counterZ0Z_24\
        );

    \I__9275\ : InMux
    port map (
            O => \N__41407\,
            I => \N__41402\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41397\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41405\,
            I => \N__41397\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__41402\,
            I => \N__41394\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__41397\,
            I => \N__41391\
        );

    \I__9270\ : Span4Mux_v
    port map (
            O => \N__41394\,
            I => \N__41388\
        );

    \I__9269\ : Span4Mux_h
    port map (
            O => \N__41391\,
            I => \N__41385\
        );

    \I__9268\ : Span4Mux_v
    port map (
            O => \N__41388\,
            I => \N__41381\
        );

    \I__9267\ : Span4Mux_v
    port map (
            O => \N__41385\,
            I => \N__41378\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41384\,
            I => \N__41375\
        );

    \I__9265\ : Odrv4
    port map (
            O => \N__41381\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__9264\ : Odrv4
    port map (
            O => \N__41378\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__41375\,
            I => \current_shift_inst.elapsed_time_ns_phase_27\
        );

    \I__9262\ : InMux
    port map (
            O => \N__41368\,
            I => \bfn_16_25_0_\
        );

    \I__9261\ : CascadeMux
    port map (
            O => \N__41365\,
            I => \N__41361\
        );

    \I__9260\ : InMux
    port map (
            O => \N__41364\,
            I => \N__41358\
        );

    \I__9259\ : InMux
    port map (
            O => \N__41361\,
            I => \N__41355\
        );

    \I__9258\ : LocalMux
    port map (
            O => \N__41358\,
            I => \N__41349\
        );

    \I__9257\ : LocalMux
    port map (
            O => \N__41355\,
            I => \N__41349\
        );

    \I__9256\ : InMux
    port map (
            O => \N__41354\,
            I => \N__41346\
        );

    \I__9255\ : Span4Mux_v
    port map (
            O => \N__41349\,
            I => \N__41343\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__41346\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__9253\ : Odrv4
    port map (
            O => \N__41343\,
            I => \current_shift_inst.timer_phase.counterZ0Z_25\
        );

    \I__9252\ : InMux
    port map (
            O => \N__41338\,
            I => \N__41333\
        );

    \I__9251\ : InMux
    port map (
            O => \N__41337\,
            I => \N__41330\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41336\,
            I => \N__41327\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__41333\,
            I => \N__41324\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__41330\,
            I => \N__41321\
        );

    \I__9247\ : LocalMux
    port map (
            O => \N__41327\,
            I => \N__41318\
        );

    \I__9246\ : Span4Mux_h
    port map (
            O => \N__41324\,
            I => \N__41315\
        );

    \I__9245\ : Span4Mux_h
    port map (
            O => \N__41321\,
            I => \N__41312\
        );

    \I__9244\ : Span12Mux_v
    port map (
            O => \N__41318\,
            I => \N__41308\
        );

    \I__9243\ : Span4Mux_v
    port map (
            O => \N__41315\,
            I => \N__41305\
        );

    \I__9242\ : Span4Mux_v
    port map (
            O => \N__41312\,
            I => \N__41302\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41311\,
            I => \N__41299\
        );

    \I__9240\ : Odrv12
    port map (
            O => \N__41308\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__9239\ : Odrv4
    port map (
            O => \N__41305\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__9238\ : Odrv4
    port map (
            O => \N__41302\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__41299\,
            I => \current_shift_inst.elapsed_time_ns_phase_28\
        );

    \I__9236\ : InMux
    port map (
            O => \N__41290\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41287\,
            I => \N__41283\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41286\,
            I => \N__41280\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__41283\,
            I => \N__41277\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__41280\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__9231\ : Odrv12
    port map (
            O => \N__41277\,
            I => \current_shift_inst.timer_phase.counterZ0Z_28\
        );

    \I__9230\ : CascadeMux
    port map (
            O => \N__41272\,
            I => \N__41267\
        );

    \I__9229\ : CascadeMux
    port map (
            O => \N__41271\,
            I => \N__41264\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41270\,
            I => \N__41261\
        );

    \I__9227\ : InMux
    port map (
            O => \N__41267\,
            I => \N__41256\
        );

    \I__9226\ : InMux
    port map (
            O => \N__41264\,
            I => \N__41256\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__41261\,
            I => \N__41251\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__41256\,
            I => \N__41251\
        );

    \I__9223\ : Odrv4
    port map (
            O => \N__41251\,
            I => \current_shift_inst.timer_phase.counterZ0Z_26\
        );

    \I__9222\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41244\
        );

    \I__9221\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41241\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__41244\,
            I => \N__41238\
        );

    \I__9219\ : LocalMux
    port map (
            O => \N__41241\,
            I => \N__41235\
        );

    \I__9218\ : Span4Mux_v
    port map (
            O => \N__41238\,
            I => \N__41232\
        );

    \I__9217\ : Span12Mux_v
    port map (
            O => \N__41235\,
            I => \N__41228\
        );

    \I__9216\ : Span4Mux_h
    port map (
            O => \N__41232\,
            I => \N__41225\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41231\,
            I => \N__41222\
        );

    \I__9214\ : Odrv12
    port map (
            O => \N__41228\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__9213\ : Odrv4
    port map (
            O => \N__41225\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__9212\ : LocalMux
    port map (
            O => \N__41222\,
            I => \current_shift_inst.elapsed_time_ns_phase_29\
        );

    \I__9211\ : InMux
    port map (
            O => \N__41215\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\
        );

    \I__9210\ : InMux
    port map (
            O => \N__41212\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\
        );

    \I__9209\ : InMux
    port map (
            O => \N__41209\,
            I => \N__41202\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41208\,
            I => \N__41202\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41207\,
            I => \N__41199\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__41202\,
            I => \N__41196\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41199\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__9204\ : Odrv12
    port map (
            O => \N__41196\,
            I => \current_shift_inst.timer_phase.counterZ0Z_12\
        );

    \I__9203\ : InMux
    port map (
            O => \N__41191\,
            I => \N__41187\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41184\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__41187\,
            I => \N__41180\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41184\,
            I => \N__41177\
        );

    \I__9199\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41174\
        );

    \I__9198\ : Span4Mux_v
    port map (
            O => \N__41180\,
            I => \N__41171\
        );

    \I__9197\ : Span4Mux_h
    port map (
            O => \N__41177\,
            I => \N__41166\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__41174\,
            I => \N__41166\
        );

    \I__9195\ : Span4Mux_v
    port map (
            O => \N__41171\,
            I => \N__41163\
        );

    \I__9194\ : Span4Mux_v
    port map (
            O => \N__41166\,
            I => \N__41160\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__41163\,
            I => \N__41156\
        );

    \I__9192\ : Span4Mux_h
    port map (
            O => \N__41160\,
            I => \N__41153\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41150\
        );

    \I__9190\ : Odrv4
    port map (
            O => \N__41156\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__9189\ : Odrv4
    port map (
            O => \N__41153\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41150\,
            I => \current_shift_inst.elapsed_time_ns_phase_15\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41143\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\
        );

    \I__9186\ : CascadeMux
    port map (
            O => \N__41140\,
            I => \N__41136\
        );

    \I__9185\ : CascadeMux
    port map (
            O => \N__41139\,
            I => \N__41133\
        );

    \I__9184\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41127\
        );

    \I__9183\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41127\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41124\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__41127\,
            I => \N__41121\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41124\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__9179\ : Odrv4
    port map (
            O => \N__41121\,
            I => \current_shift_inst.timer_phase.counterZ0Z_13\
        );

    \I__9178\ : CascadeMux
    port map (
            O => \N__41116\,
            I => \N__41112\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41115\,
            I => \N__41108\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41112\,
            I => \N__41105\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41111\,
            I => \N__41102\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41108\,
            I => \N__41099\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__41105\,
            I => \N__41094\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__41102\,
            I => \N__41094\
        );

    \I__9171\ : Span4Mux_h
    port map (
            O => \N__41099\,
            I => \N__41091\
        );

    \I__9170\ : Span12Mux_h
    port map (
            O => \N__41094\,
            I => \N__41087\
        );

    \I__9169\ : Span4Mux_v
    port map (
            O => \N__41091\,
            I => \N__41084\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41090\,
            I => \N__41081\
        );

    \I__9167\ : Odrv12
    port map (
            O => \N__41087\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__9166\ : Odrv4
    port map (
            O => \N__41084\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__9165\ : LocalMux
    port map (
            O => \N__41081\,
            I => \current_shift_inst.elapsed_time_ns_phase_16\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41074\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\
        );

    \I__9163\ : CascadeMux
    port map (
            O => \N__41071\,
            I => \N__41067\
        );

    \I__9162\ : CascadeMux
    port map (
            O => \N__41070\,
            I => \N__41064\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41067\,
            I => \N__41058\
        );

    \I__9160\ : InMux
    port map (
            O => \N__41064\,
            I => \N__41058\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41063\,
            I => \N__41055\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41058\,
            I => \N__41052\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41055\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__9156\ : Odrv12
    port map (
            O => \N__41052\,
            I => \current_shift_inst.timer_phase.counterZ0Z_14\
        );

    \I__9155\ : InMux
    port map (
            O => \N__41047\,
            I => \N__41044\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41044\,
            I => \N__41040\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41043\,
            I => \N__41037\
        );

    \I__9152\ : Span4Mux_h
    port map (
            O => \N__41040\,
            I => \N__41031\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__41037\,
            I => \N__41031\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41036\,
            I => \N__41028\
        );

    \I__9149\ : Span4Mux_h
    port map (
            O => \N__41031\,
            I => \N__41025\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41028\,
            I => \N__41022\
        );

    \I__9147\ : Span4Mux_v
    port map (
            O => \N__41025\,
            I => \N__41018\
        );

    \I__9146\ : Span12Mux_h
    port map (
            O => \N__41022\,
            I => \N__41015\
        );

    \I__9145\ : InMux
    port map (
            O => \N__41021\,
            I => \N__41012\
        );

    \I__9144\ : Odrv4
    port map (
            O => \N__41018\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__9143\ : Odrv12
    port map (
            O => \N__41015\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__41012\,
            I => \current_shift_inst.elapsed_time_ns_phase_17\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41005\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41002\,
            I => \N__40995\
        );

    \I__9139\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40995\
        );

    \I__9138\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40992\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__40995\,
            I => \N__40989\
        );

    \I__9136\ : LocalMux
    port map (
            O => \N__40992\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__9135\ : Odrv12
    port map (
            O => \N__40989\,
            I => \current_shift_inst.timer_phase.counterZ0Z_15\
        );

    \I__9134\ : InMux
    port map (
            O => \N__40984\,
            I => \N__40979\
        );

    \I__9133\ : InMux
    port map (
            O => \N__40983\,
            I => \N__40974\
        );

    \I__9132\ : InMux
    port map (
            O => \N__40982\,
            I => \N__40974\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40971\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__40974\,
            I => \N__40968\
        );

    \I__9129\ : Span4Mux_h
    port map (
            O => \N__40971\,
            I => \N__40965\
        );

    \I__9128\ : Span4Mux_h
    port map (
            O => \N__40968\,
            I => \N__40962\
        );

    \I__9127\ : Span4Mux_v
    port map (
            O => \N__40965\,
            I => \N__40959\
        );

    \I__9126\ : Span4Mux_v
    port map (
            O => \N__40962\,
            I => \N__40955\
        );

    \I__9125\ : Span4Mux_h
    port map (
            O => \N__40959\,
            I => \N__40952\
        );

    \I__9124\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40949\
        );

    \I__9123\ : Odrv4
    port map (
            O => \N__40955\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__40952\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__40949\,
            I => \current_shift_inst.elapsed_time_ns_phase_18\
        );

    \I__9120\ : InMux
    port map (
            O => \N__40942\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\
        );

    \I__9119\ : InMux
    port map (
            O => \N__40939\,
            I => \N__40935\
        );

    \I__9118\ : InMux
    port map (
            O => \N__40938\,
            I => \N__40932\
        );

    \I__9117\ : LocalMux
    port map (
            O => \N__40935\,
            I => \N__40929\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__40932\,
            I => \N__40923\
        );

    \I__9115\ : Span4Mux_v
    port map (
            O => \N__40929\,
            I => \N__40923\
        );

    \I__9114\ : InMux
    port map (
            O => \N__40928\,
            I => \N__40920\
        );

    \I__9113\ : Span4Mux_h
    port map (
            O => \N__40923\,
            I => \N__40917\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__40920\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__9111\ : Odrv4
    port map (
            O => \N__40917\,
            I => \current_shift_inst.timer_phase.counterZ0Z_16\
        );

    \I__9110\ : InMux
    port map (
            O => \N__40912\,
            I => \N__40906\
        );

    \I__9109\ : InMux
    port map (
            O => \N__40911\,
            I => \N__40906\
        );

    \I__9108\ : LocalMux
    port map (
            O => \N__40906\,
            I => \N__40902\
        );

    \I__9107\ : InMux
    port map (
            O => \N__40905\,
            I => \N__40899\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__40902\,
            I => \N__40894\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__40899\,
            I => \N__40894\
        );

    \I__9104\ : Span4Mux_v
    port map (
            O => \N__40894\,
            I => \N__40891\
        );

    \I__9103\ : Span4Mux_v
    port map (
            O => \N__40891\,
            I => \N__40888\
        );

    \I__9102\ : Span4Mux_h
    port map (
            O => \N__40888\,
            I => \N__40884\
        );

    \I__9101\ : InMux
    port map (
            O => \N__40887\,
            I => \N__40881\
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__40884\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__40881\,
            I => \current_shift_inst.elapsed_time_ns_phase_19\
        );

    \I__9098\ : InMux
    port map (
            O => \N__40876\,
            I => \bfn_16_24_0_\
        );

    \I__9097\ : CascadeMux
    port map (
            O => \N__40873\,
            I => \N__40870\
        );

    \I__9096\ : InMux
    port map (
            O => \N__40870\,
            I => \N__40867\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__40867\,
            I => \N__40863\
        );

    \I__9094\ : InMux
    port map (
            O => \N__40866\,
            I => \N__40859\
        );

    \I__9093\ : Span4Mux_v
    port map (
            O => \N__40863\,
            I => \N__40856\
        );

    \I__9092\ : InMux
    port map (
            O => \N__40862\,
            I => \N__40853\
        );

    \I__9091\ : LocalMux
    port map (
            O => \N__40859\,
            I => \N__40848\
        );

    \I__9090\ : Span4Mux_h
    port map (
            O => \N__40856\,
            I => \N__40848\
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__40853\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__9088\ : Odrv4
    port map (
            O => \N__40848\,
            I => \current_shift_inst.timer_phase.counterZ0Z_17\
        );

    \I__9087\ : InMux
    port map (
            O => \N__40843\,
            I => \N__40839\
        );

    \I__9086\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40835\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__40839\,
            I => \N__40832\
        );

    \I__9084\ : InMux
    port map (
            O => \N__40838\,
            I => \N__40829\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__40835\,
            I => \N__40826\
        );

    \I__9082\ : Span4Mux_h
    port map (
            O => \N__40832\,
            I => \N__40821\
        );

    \I__9081\ : LocalMux
    port map (
            O => \N__40829\,
            I => \N__40821\
        );

    \I__9080\ : Sp12to4
    port map (
            O => \N__40826\,
            I => \N__40818\
        );

    \I__9079\ : Span4Mux_h
    port map (
            O => \N__40821\,
            I => \N__40815\
        );

    \I__9078\ : Span12Mux_v
    port map (
            O => \N__40818\,
            I => \N__40811\
        );

    \I__9077\ : Span4Mux_v
    port map (
            O => \N__40815\,
            I => \N__40808\
        );

    \I__9076\ : InMux
    port map (
            O => \N__40814\,
            I => \N__40805\
        );

    \I__9075\ : Odrv12
    port map (
            O => \N__40811\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__9074\ : Odrv4
    port map (
            O => \N__40808\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__9073\ : LocalMux
    port map (
            O => \N__40805\,
            I => \current_shift_inst.elapsed_time_ns_phase_20\
        );

    \I__9072\ : InMux
    port map (
            O => \N__40798\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\
        );

    \I__9071\ : CascadeMux
    port map (
            O => \N__40795\,
            I => \N__40790\
        );

    \I__9070\ : InMux
    port map (
            O => \N__40794\,
            I => \N__40787\
        );

    \I__9069\ : InMux
    port map (
            O => \N__40793\,
            I => \N__40784\
        );

    \I__9068\ : InMux
    port map (
            O => \N__40790\,
            I => \N__40781\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__40787\,
            I => \N__40774\
        );

    \I__9066\ : LocalMux
    port map (
            O => \N__40784\,
            I => \N__40774\
        );

    \I__9065\ : LocalMux
    port map (
            O => \N__40781\,
            I => \N__40774\
        );

    \I__9064\ : Odrv4
    port map (
            O => \N__40774\,
            I => \current_shift_inst.timer_phase.counterZ0Z_18\
        );

    \I__9063\ : InMux
    port map (
            O => \N__40771\,
            I => \N__40765\
        );

    \I__9062\ : InMux
    port map (
            O => \N__40770\,
            I => \N__40765\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__40765\,
            I => \N__40761\
        );

    \I__9060\ : InMux
    port map (
            O => \N__40764\,
            I => \N__40758\
        );

    \I__9059\ : Span4Mux_h
    port map (
            O => \N__40761\,
            I => \N__40755\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__40758\,
            I => \N__40752\
        );

    \I__9057\ : Span4Mux_v
    port map (
            O => \N__40755\,
            I => \N__40749\
        );

    \I__9056\ : Span12Mux_h
    port map (
            O => \N__40752\,
            I => \N__40745\
        );

    \I__9055\ : Span4Mux_h
    port map (
            O => \N__40749\,
            I => \N__40742\
        );

    \I__9054\ : InMux
    port map (
            O => \N__40748\,
            I => \N__40739\
        );

    \I__9053\ : Odrv12
    port map (
            O => \N__40745\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__9052\ : Odrv4
    port map (
            O => \N__40742\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__40739\,
            I => \current_shift_inst.elapsed_time_ns_phase_21\
        );

    \I__9050\ : InMux
    port map (
            O => \N__40732\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\
        );

    \I__9049\ : CascadeMux
    port map (
            O => \N__40729\,
            I => \N__40725\
        );

    \I__9048\ : CascadeMux
    port map (
            O => \N__40728\,
            I => \N__40722\
        );

    \I__9047\ : InMux
    port map (
            O => \N__40725\,
            I => \N__40716\
        );

    \I__9046\ : InMux
    port map (
            O => \N__40722\,
            I => \N__40716\
        );

    \I__9045\ : InMux
    port map (
            O => \N__40721\,
            I => \N__40713\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__40716\,
            I => \N__40710\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__40713\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__40710\,
            I => \current_shift_inst.timer_phase.counterZ0Z_4\
        );

    \I__9041\ : CascadeMux
    port map (
            O => \N__40705\,
            I => \N__40702\
        );

    \I__9040\ : InMux
    port map (
            O => \N__40702\,
            I => \N__40698\
        );

    \I__9039\ : CascadeMux
    port map (
            O => \N__40701\,
            I => \N__40694\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__40698\,
            I => \N__40691\
        );

    \I__9037\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40686\
        );

    \I__9036\ : InMux
    port map (
            O => \N__40694\,
            I => \N__40686\
        );

    \I__9035\ : Span4Mux_v
    port map (
            O => \N__40691\,
            I => \N__40683\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__40686\,
            I => \N__40680\
        );

    \I__9033\ : Span4Mux_h
    port map (
            O => \N__40683\,
            I => \N__40676\
        );

    \I__9032\ : Sp12to4
    port map (
            O => \N__40680\,
            I => \N__40673\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40679\,
            I => \N__40670\
        );

    \I__9030\ : Odrv4
    port map (
            O => \N__40676\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__9029\ : Odrv12
    port map (
            O => \N__40673\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__40670\,
            I => \current_shift_inst.elapsed_time_ns_phase_7\
        );

    \I__9027\ : InMux
    port map (
            O => \N__40663\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__40660\,
            I => \N__40656\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__40659\,
            I => \N__40653\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40656\,
            I => \N__40647\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40647\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40652\,
            I => \N__40644\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__40647\,
            I => \N__40641\
        );

    \I__9020\ : LocalMux
    port map (
            O => \N__40644\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__9019\ : Odrv4
    port map (
            O => \N__40641\,
            I => \current_shift_inst.timer_phase.counterZ0Z_5\
        );

    \I__9018\ : CascadeMux
    port map (
            O => \N__40636\,
            I => \N__40633\
        );

    \I__9017\ : InMux
    port map (
            O => \N__40633\,
            I => \N__40629\
        );

    \I__9016\ : InMux
    port map (
            O => \N__40632\,
            I => \N__40625\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__40629\,
            I => \N__40622\
        );

    \I__9014\ : InMux
    port map (
            O => \N__40628\,
            I => \N__40619\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__40625\,
            I => \N__40616\
        );

    \I__9012\ : Span4Mux_v
    port map (
            O => \N__40622\,
            I => \N__40613\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__40619\,
            I => \N__40610\
        );

    \I__9010\ : Span4Mux_h
    port map (
            O => \N__40616\,
            I => \N__40607\
        );

    \I__9009\ : Span4Mux_h
    port map (
            O => \N__40613\,
            I => \N__40603\
        );

    \I__9008\ : Span4Mux_h
    port map (
            O => \N__40610\,
            I => \N__40600\
        );

    \I__9007\ : Span4Mux_v
    port map (
            O => \N__40607\,
            I => \N__40597\
        );

    \I__9006\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40594\
        );

    \I__9005\ : Odrv4
    port map (
            O => \N__40603\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__9004\ : Odrv4
    port map (
            O => \N__40600\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__9003\ : Odrv4
    port map (
            O => \N__40597\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__9002\ : LocalMux
    port map (
            O => \N__40594\,
            I => \current_shift_inst.elapsed_time_ns_phase_8\
        );

    \I__9001\ : InMux
    port map (
            O => \N__40585\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\
        );

    \I__9000\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40575\
        );

    \I__8999\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40575\
        );

    \I__8998\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40572\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__40575\,
            I => \N__40569\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__40572\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__8995\ : Odrv12
    port map (
            O => \N__40569\,
            I => \current_shift_inst.timer_phase.counterZ0Z_6\
        );

    \I__8994\ : InMux
    port map (
            O => \N__40564\,
            I => \N__40557\
        );

    \I__8993\ : InMux
    port map (
            O => \N__40563\,
            I => \N__40557\
        );

    \I__8992\ : InMux
    port map (
            O => \N__40562\,
            I => \N__40554\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__40557\,
            I => \N__40551\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__40554\,
            I => \N__40548\
        );

    \I__8989\ : Span4Mux_h
    port map (
            O => \N__40551\,
            I => \N__40545\
        );

    \I__8988\ : Span4Mux_h
    port map (
            O => \N__40548\,
            I => \N__40542\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__40545\,
            I => \N__40538\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__40542\,
            I => \N__40535\
        );

    \I__8985\ : InMux
    port map (
            O => \N__40541\,
            I => \N__40532\
        );

    \I__8984\ : Odrv4
    port map (
            O => \N__40538\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__8983\ : Odrv4
    port map (
            O => \N__40535\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__40532\,
            I => \current_shift_inst.elapsed_time_ns_phase_9\
        );

    \I__8981\ : InMux
    port map (
            O => \N__40525\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\
        );

    \I__8980\ : InMux
    port map (
            O => \N__40522\,
            I => \N__40515\
        );

    \I__8979\ : InMux
    port map (
            O => \N__40521\,
            I => \N__40515\
        );

    \I__8978\ : InMux
    port map (
            O => \N__40520\,
            I => \N__40512\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__40515\,
            I => \N__40509\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__40512\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__8975\ : Odrv12
    port map (
            O => \N__40509\,
            I => \current_shift_inst.timer_phase.counterZ0Z_7\
        );

    \I__8974\ : InMux
    port map (
            O => \N__40504\,
            I => \N__40499\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40503\,
            I => \N__40496\
        );

    \I__8972\ : InMux
    port map (
            O => \N__40502\,
            I => \N__40493\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__40499\,
            I => \N__40490\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__40496\,
            I => \N__40487\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__40493\,
            I => \N__40484\
        );

    \I__8968\ : Span4Mux_h
    port map (
            O => \N__40490\,
            I => \N__40481\
        );

    \I__8967\ : Span4Mux_h
    port map (
            O => \N__40487\,
            I => \N__40478\
        );

    \I__8966\ : Span4Mux_v
    port map (
            O => \N__40484\,
            I => \N__40473\
        );

    \I__8965\ : Span4Mux_v
    port map (
            O => \N__40481\,
            I => \N__40473\
        );

    \I__8964\ : Span4Mux_h
    port map (
            O => \N__40478\,
            I => \N__40469\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__40473\,
            I => \N__40466\
        );

    \I__8962\ : InMux
    port map (
            O => \N__40472\,
            I => \N__40463\
        );

    \I__8961\ : Odrv4
    port map (
            O => \N__40469\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__8960\ : Odrv4
    port map (
            O => \N__40466\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__40463\,
            I => \current_shift_inst.elapsed_time_ns_phase_10\
        );

    \I__8958\ : InMux
    port map (
            O => \N__40456\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\
        );

    \I__8957\ : CascadeMux
    port map (
            O => \N__40453\,
            I => \N__40450\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40447\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__40447\,
            I => \N__40443\
        );

    \I__8954\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40439\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__40443\,
            I => \N__40436\
        );

    \I__8952\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40433\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__40439\,
            I => \N__40428\
        );

    \I__8950\ : Span4Mux_h
    port map (
            O => \N__40436\,
            I => \N__40428\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__40433\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__8948\ : Odrv4
    port map (
            O => \N__40428\,
            I => \current_shift_inst.timer_phase.counterZ0Z_8\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__40423\,
            I => \N__40420\
        );

    \I__8946\ : InMux
    port map (
            O => \N__40420\,
            I => \N__40416\
        );

    \I__8945\ : InMux
    port map (
            O => \N__40419\,
            I => \N__40413\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__40416\,
            I => \N__40409\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__40413\,
            I => \N__40406\
        );

    \I__8942\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40403\
        );

    \I__8941\ : Span4Mux_h
    port map (
            O => \N__40409\,
            I => \N__40400\
        );

    \I__8940\ : Span4Mux_h
    port map (
            O => \N__40406\,
            I => \N__40397\
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__40403\,
            I => \N__40394\
        );

    \I__8938\ : Span4Mux_v
    port map (
            O => \N__40400\,
            I => \N__40390\
        );

    \I__8937\ : Span4Mux_h
    port map (
            O => \N__40397\,
            I => \N__40387\
        );

    \I__8936\ : Span12Mux_h
    port map (
            O => \N__40394\,
            I => \N__40384\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40393\,
            I => \N__40381\
        );

    \I__8934\ : Odrv4
    port map (
            O => \N__40390\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__8933\ : Odrv4
    port map (
            O => \N__40387\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__8932\ : Odrv12
    port map (
            O => \N__40384\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__40381\,
            I => \current_shift_inst.elapsed_time_ns_phase_11\
        );

    \I__8930\ : InMux
    port map (
            O => \N__40372\,
            I => \bfn_16_23_0_\
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__40369\,
            I => \N__40365\
        );

    \I__8928\ : InMux
    port map (
            O => \N__40368\,
            I => \N__40362\
        );

    \I__8927\ : InMux
    port map (
            O => \N__40365\,
            I => \N__40359\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__40362\,
            I => \N__40353\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__40359\,
            I => \N__40353\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40358\,
            I => \N__40350\
        );

    \I__8923\ : Span4Mux_v
    port map (
            O => \N__40353\,
            I => \N__40347\
        );

    \I__8922\ : LocalMux
    port map (
            O => \N__40350\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__8921\ : Odrv4
    port map (
            O => \N__40347\,
            I => \current_shift_inst.timer_phase.counterZ0Z_9\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40342\,
            I => \N__40337\
        );

    \I__8919\ : InMux
    port map (
            O => \N__40341\,
            I => \N__40332\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40340\,
            I => \N__40332\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__40337\,
            I => \N__40329\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__40332\,
            I => \N__40326\
        );

    \I__8915\ : Span4Mux_h
    port map (
            O => \N__40329\,
            I => \N__40323\
        );

    \I__8914\ : Span4Mux_h
    port map (
            O => \N__40326\,
            I => \N__40320\
        );

    \I__8913\ : Span4Mux_h
    port map (
            O => \N__40323\,
            I => \N__40316\
        );

    \I__8912\ : Span4Mux_v
    port map (
            O => \N__40320\,
            I => \N__40313\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40319\,
            I => \N__40310\
        );

    \I__8910\ : Odrv4
    port map (
            O => \N__40316\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__8909\ : Odrv4
    port map (
            O => \N__40313\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__40310\,
            I => \current_shift_inst.elapsed_time_ns_phase_12\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40303\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\
        );

    \I__8906\ : CascadeMux
    port map (
            O => \N__40300\,
            I => \N__40295\
        );

    \I__8905\ : CascadeMux
    port map (
            O => \N__40299\,
            I => \N__40292\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40298\,
            I => \N__40289\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40295\,
            I => \N__40284\
        );

    \I__8902\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40284\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__40289\,
            I => \N__40279\
        );

    \I__8900\ : LocalMux
    port map (
            O => \N__40284\,
            I => \N__40279\
        );

    \I__8899\ : Odrv4
    port map (
            O => \N__40279\,
            I => \current_shift_inst.timer_phase.counterZ0Z_10\
        );

    \I__8898\ : CascadeMux
    port map (
            O => \N__40276\,
            I => \N__40273\
        );

    \I__8897\ : InMux
    port map (
            O => \N__40273\,
            I => \N__40270\
        );

    \I__8896\ : LocalMux
    port map (
            O => \N__40270\,
            I => \N__40266\
        );

    \I__8895\ : InMux
    port map (
            O => \N__40269\,
            I => \N__40262\
        );

    \I__8894\ : Span4Mux_h
    port map (
            O => \N__40266\,
            I => \N__40259\
        );

    \I__8893\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40256\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__40262\,
            I => \N__40253\
        );

    \I__8891\ : Span4Mux_h
    port map (
            O => \N__40259\,
            I => \N__40250\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__40256\,
            I => \N__40247\
        );

    \I__8889\ : Span4Mux_h
    port map (
            O => \N__40253\,
            I => \N__40244\
        );

    \I__8888\ : Sp12to4
    port map (
            O => \N__40250\,
            I => \N__40240\
        );

    \I__8887\ : Span12Mux_h
    port map (
            O => \N__40247\,
            I => \N__40237\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__40244\,
            I => \N__40234\
        );

    \I__8885\ : InMux
    port map (
            O => \N__40243\,
            I => \N__40231\
        );

    \I__8884\ : Odrv12
    port map (
            O => \N__40240\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__8883\ : Odrv12
    port map (
            O => \N__40237\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__8882\ : Odrv4
    port map (
            O => \N__40234\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__40231\,
            I => \current_shift_inst.elapsed_time_ns_phase_13\
        );

    \I__8880\ : InMux
    port map (
            O => \N__40222\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\
        );

    \I__8879\ : CascadeMux
    port map (
            O => \N__40219\,
            I => \N__40214\
        );

    \I__8878\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40211\
        );

    \I__8877\ : InMux
    port map (
            O => \N__40217\,
            I => \N__40208\
        );

    \I__8876\ : InMux
    port map (
            O => \N__40214\,
            I => \N__40205\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__40211\,
            I => \N__40198\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__40208\,
            I => \N__40198\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40205\,
            I => \N__40198\
        );

    \I__8872\ : Odrv4
    port map (
            O => \N__40198\,
            I => \current_shift_inst.timer_phase.counterZ0Z_11\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40195\,
            I => \N__40190\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40194\,
            I => \N__40187\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40193\,
            I => \N__40184\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40190\,
            I => \N__40181\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__40187\,
            I => \N__40178\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__40184\,
            I => \N__40175\
        );

    \I__8865\ : Span4Mux_h
    port map (
            O => \N__40181\,
            I => \N__40170\
        );

    \I__8864\ : Span4Mux_v
    port map (
            O => \N__40178\,
            I => \N__40170\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__40175\,
            I => \N__40167\
        );

    \I__8862\ : Span4Mux_v
    port map (
            O => \N__40170\,
            I => \N__40164\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__40167\,
            I => \N__40160\
        );

    \I__8860\ : Span4Mux_h
    port map (
            O => \N__40164\,
            I => \N__40157\
        );

    \I__8859\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40154\
        );

    \I__8858\ : Odrv4
    port map (
            O => \N__40160\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__8857\ : Odrv4
    port map (
            O => \N__40157\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__8856\ : LocalMux
    port map (
            O => \N__40154\,
            I => \current_shift_inst.elapsed_time_ns_phase_14\
        );

    \I__8855\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40144\
        );

    \I__8854\ : LocalMux
    port map (
            O => \N__40144\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5\
        );

    \I__8853\ : CascadeMux
    port map (
            O => \N__40141\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4_cascade_\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40138\,
            I => \N__40135\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__8850\ : Odrv4
    port map (
            O => \N__40132\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6\
        );

    \I__8849\ : InMux
    port map (
            O => \N__40129\,
            I => \N__40126\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__40126\,
            I => \N__40122\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40125\,
            I => \N__40119\
        );

    \I__8846\ : Span4Mux_h
    port map (
            O => \N__40122\,
            I => \N__40115\
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40119\,
            I => \N__40112\
        );

    \I__8844\ : InMux
    port map (
            O => \N__40118\,
            I => \N__40109\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__40115\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__40112\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__8841\ : LocalMux
    port map (
            O => \N__40109\,
            I => \current_shift_inst.timer_phase.counterZ0Z_0\
        );

    \I__8840\ : InMux
    port map (
            O => \N__40102\,
            I => \N__40096\
        );

    \I__8839\ : InMux
    port map (
            O => \N__40101\,
            I => \N__40096\
        );

    \I__8838\ : LocalMux
    port map (
            O => \N__40096\,
            I => \N__40092\
        );

    \I__8837\ : InMux
    port map (
            O => \N__40095\,
            I => \N__40089\
        );

    \I__8836\ : Odrv4
    port map (
            O => \N__40092\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__40089\,
            I => \current_shift_inst.elapsed_time_ns_phase_3\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40084\,
            I => \N__40079\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40083\,
            I => \N__40076\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40082\,
            I => \N__40073\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40079\,
            I => \N__40070\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__40076\,
            I => \N__40065\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40073\,
            I => \N__40065\
        );

    \I__8828\ : Odrv4
    port map (
            O => \N__40070\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__8827\ : Odrv4
    port map (
            O => \N__40065\,
            I => \current_shift_inst.timer_phase.counterZ0Z_1\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40060\,
            I => \N__40053\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40053\
        );

    \I__8824\ : InMux
    port map (
            O => \N__40058\,
            I => \N__40050\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40053\,
            I => \N__40047\
        );

    \I__8822\ : LocalMux
    port map (
            O => \N__40050\,
            I => \N__40044\
        );

    \I__8821\ : Span4Mux_h
    port map (
            O => \N__40047\,
            I => \N__40041\
        );

    \I__8820\ : Span4Mux_h
    port map (
            O => \N__40044\,
            I => \N__40038\
        );

    \I__8819\ : Span4Mux_h
    port map (
            O => \N__40041\,
            I => \N__40034\
        );

    \I__8818\ : Span4Mux_h
    port map (
            O => \N__40038\,
            I => \N__40031\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40037\,
            I => \N__40028\
        );

    \I__8816\ : Odrv4
    port map (
            O => \N__40034\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__8815\ : Odrv4
    port map (
            O => \N__40031\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40028\,
            I => \current_shift_inst.elapsed_time_ns_phase_4\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40021\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\
        );

    \I__8812\ : CascadeMux
    port map (
            O => \N__40018\,
            I => \N__40013\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40017\,
            I => \N__40010\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40016\,
            I => \N__40007\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40013\,
            I => \N__40004\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__40010\,
            I => \N__39997\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__40007\,
            I => \N__39997\
        );

    \I__8806\ : LocalMux
    port map (
            O => \N__40004\,
            I => \N__39997\
        );

    \I__8805\ : Odrv4
    port map (
            O => \N__39997\,
            I => \current_shift_inst.timer_phase.counterZ0Z_2\
        );

    \I__8804\ : InMux
    port map (
            O => \N__39994\,
            I => \N__39991\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__39991\,
            I => \N__39986\
        );

    \I__8802\ : InMux
    port map (
            O => \N__39990\,
            I => \N__39983\
        );

    \I__8801\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39980\
        );

    \I__8800\ : Span4Mux_v
    port map (
            O => \N__39986\,
            I => \N__39975\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__39983\,
            I => \N__39975\
        );

    \I__8798\ : LocalMux
    port map (
            O => \N__39980\,
            I => \N__39972\
        );

    \I__8797\ : Sp12to4
    port map (
            O => \N__39975\,
            I => \N__39966\
        );

    \I__8796\ : Span12Mux_v
    port map (
            O => \N__39972\,
            I => \N__39966\
        );

    \I__8795\ : InMux
    port map (
            O => \N__39971\,
            I => \N__39963\
        );

    \I__8794\ : Odrv12
    port map (
            O => \N__39966\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__39963\,
            I => \current_shift_inst.elapsed_time_ns_phase_5\
        );

    \I__8792\ : InMux
    port map (
            O => \N__39958\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\
        );

    \I__8791\ : CascadeMux
    port map (
            O => \N__39955\,
            I => \N__39950\
        );

    \I__8790\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39947\
        );

    \I__8789\ : InMux
    port map (
            O => \N__39953\,
            I => \N__39944\
        );

    \I__8788\ : InMux
    port map (
            O => \N__39950\,
            I => \N__39941\
        );

    \I__8787\ : LocalMux
    port map (
            O => \N__39947\,
            I => \N__39934\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__39944\,
            I => \N__39934\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__39941\,
            I => \N__39934\
        );

    \I__8784\ : Odrv4
    port map (
            O => \N__39934\,
            I => \current_shift_inst.timer_phase.counterZ0Z_3\
        );

    \I__8783\ : InMux
    port map (
            O => \N__39931\,
            I => \N__39926\
        );

    \I__8782\ : InMux
    port map (
            O => \N__39930\,
            I => \N__39921\
        );

    \I__8781\ : InMux
    port map (
            O => \N__39929\,
            I => \N__39921\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__39926\,
            I => \N__39918\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__39921\,
            I => \N__39914\
        );

    \I__8778\ : Span4Mux_h
    port map (
            O => \N__39918\,
            I => \N__39911\
        );

    \I__8777\ : InMux
    port map (
            O => \N__39917\,
            I => \N__39908\
        );

    \I__8776\ : Odrv12
    port map (
            O => \N__39914\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__8775\ : Odrv4
    port map (
            O => \N__39911\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__39908\,
            I => \current_shift_inst.elapsed_time_ns_phase_6\
        );

    \I__8773\ : InMux
    port map (
            O => \N__39901\,
            I => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\
        );

    \I__8772\ : InMux
    port map (
            O => \N__39898\,
            I => \N__39895\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__39895\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\
        );

    \I__8770\ : InMux
    port map (
            O => \N__39892\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__8769\ : InMux
    port map (
            O => \N__39889\,
            I => \N__39886\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__39886\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\
        );

    \I__8767\ : InMux
    port map (
            O => \N__39883\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__8766\ : CEMux
    port map (
            O => \N__39880\,
            I => \N__39862\
        );

    \I__8765\ : CEMux
    port map (
            O => \N__39879\,
            I => \N__39862\
        );

    \I__8764\ : CEMux
    port map (
            O => \N__39878\,
            I => \N__39862\
        );

    \I__8763\ : CEMux
    port map (
            O => \N__39877\,
            I => \N__39862\
        );

    \I__8762\ : CEMux
    port map (
            O => \N__39876\,
            I => \N__39862\
        );

    \I__8761\ : CEMux
    port map (
            O => \N__39875\,
            I => \N__39862\
        );

    \I__8760\ : GlobalMux
    port map (
            O => \N__39862\,
            I => \N__39859\
        );

    \I__8759\ : gio2CtrlBuf
    port map (
            O => \N__39859\,
            I => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \I__8758\ : InMux
    port map (
            O => \N__39856\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__8757\ : InMux
    port map (
            O => \N__39853\,
            I => \N__39850\
        );

    \I__8756\ : LocalMux
    port map (
            O => \N__39850\,
            I => \N__39846\
        );

    \I__8755\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39843\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__39846\,
            I => \N__39838\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__39843\,
            I => \N__39838\
        );

    \I__8752\ : Span4Mux_v
    port map (
            O => \N__39838\,
            I => \N__39835\
        );

    \I__8751\ : Odrv4
    port map (
            O => \N__39835\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__8750\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39828\
        );

    \I__8749\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39825\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__39828\,
            I => \N__39821\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__39825\,
            I => \N__39818\
        );

    \I__8746\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39815\
        );

    \I__8745\ : Span4Mux_v
    port map (
            O => \N__39821\,
            I => \N__39811\
        );

    \I__8744\ : Span12Mux_v
    port map (
            O => \N__39818\,
            I => \N__39806\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__39815\,
            I => \N__39806\
        );

    \I__8742\ : InMux
    port map (
            O => \N__39814\,
            I => \N__39803\
        );

    \I__8741\ : Span4Mux_h
    port map (
            O => \N__39811\,
            I => \N__39800\
        );

    \I__8740\ : Span12Mux_v
    port map (
            O => \N__39806\,
            I => \N__39797\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__39803\,
            I => \N__39794\
        );

    \I__8738\ : Odrv4
    port map (
            O => \N__39800\,
            I => measured_delay_tr_18
        );

    \I__8737\ : Odrv12
    port map (
            O => \N__39797\,
            I => measured_delay_tr_18
        );

    \I__8736\ : Odrv4
    port map (
            O => \N__39794\,
            I => measured_delay_tr_18
        );

    \I__8735\ : InMux
    port map (
            O => \N__39787\,
            I => \N__39783\
        );

    \I__8734\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39779\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__39783\,
            I => \N__39776\
        );

    \I__8732\ : InMux
    port map (
            O => \N__39782\,
            I => \N__39773\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__39779\,
            I => \N__39770\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__39776\,
            I => \N__39767\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__39773\,
            I => \N__39764\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__39770\,
            I => \N__39760\
        );

    \I__8727\ : Span4Mux_v
    port map (
            O => \N__39767\,
            I => \N__39755\
        );

    \I__8726\ : Span4Mux_v
    port map (
            O => \N__39764\,
            I => \N__39755\
        );

    \I__8725\ : InMux
    port map (
            O => \N__39763\,
            I => \N__39752\
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__39760\,
            I => measured_delay_tr_17
        );

    \I__8723\ : Odrv4
    port map (
            O => \N__39755\,
            I => measured_delay_tr_17
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__39752\,
            I => measured_delay_tr_17
        );

    \I__8721\ : CascadeMux
    port map (
            O => \N__39745\,
            I => \N__39742\
        );

    \I__8720\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39737\
        );

    \I__8719\ : InMux
    port map (
            O => \N__39741\,
            I => \N__39733\
        );

    \I__8718\ : InMux
    port map (
            O => \N__39740\,
            I => \N__39730\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__39737\,
            I => \N__39727\
        );

    \I__8716\ : CascadeMux
    port map (
            O => \N__39736\,
            I => \N__39724\
        );

    \I__8715\ : LocalMux
    port map (
            O => \N__39733\,
            I => \N__39721\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__39730\,
            I => \N__39718\
        );

    \I__8713\ : Span4Mux_v
    port map (
            O => \N__39727\,
            I => \N__39715\
        );

    \I__8712\ : InMux
    port map (
            O => \N__39724\,
            I => \N__39712\
        );

    \I__8711\ : Span12Mux_h
    port map (
            O => \N__39721\,
            I => \N__39709\
        );

    \I__8710\ : Span4Mux_v
    port map (
            O => \N__39718\,
            I => \N__39706\
        );

    \I__8709\ : Span4Mux_h
    port map (
            O => \N__39715\,
            I => \N__39701\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__39712\,
            I => \N__39701\
        );

    \I__8707\ : Odrv12
    port map (
            O => \N__39709\,
            I => measured_delay_tr_19
        );

    \I__8706\ : Odrv4
    port map (
            O => \N__39706\,
            I => measured_delay_tr_19
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__39701\,
            I => measured_delay_tr_19
        );

    \I__8704\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39691\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__39691\,
            I => \N__39687\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39690\,
            I => \N__39684\
        );

    \I__8701\ : Span4Mux_h
    port map (
            O => \N__39687\,
            I => \N__39680\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__39684\,
            I => \N__39677\
        );

    \I__8699\ : CascadeMux
    port map (
            O => \N__39683\,
            I => \N__39674\
        );

    \I__8698\ : Span4Mux_v
    port map (
            O => \N__39680\,
            I => \N__39670\
        );

    \I__8697\ : Span4Mux_h
    port map (
            O => \N__39677\,
            I => \N__39667\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39674\,
            I => \N__39663\
        );

    \I__8695\ : InMux
    port map (
            O => \N__39673\,
            I => \N__39660\
        );

    \I__8694\ : Span4Mux_v
    port map (
            O => \N__39670\,
            I => \N__39655\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__39667\,
            I => \N__39655\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39652\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__39663\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__39660\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8689\ : Odrv4
    port map (
            O => \N__39655\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8688\ : LocalMux
    port map (
            O => \N__39652\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__8687\ : InMux
    port map (
            O => \N__39643\,
            I => \N__39639\
        );

    \I__8686\ : InMux
    port map (
            O => \N__39642\,
            I => \N__39636\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39632\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39628\
        );

    \I__8683\ : InMux
    port map (
            O => \N__39635\,
            I => \N__39625\
        );

    \I__8682\ : Sp12to4
    port map (
            O => \N__39632\,
            I => \N__39622\
        );

    \I__8681\ : InMux
    port map (
            O => \N__39631\,
            I => \N__39619\
        );

    \I__8680\ : Span12Mux_v
    port map (
            O => \N__39628\,
            I => \N__39616\
        );

    \I__8679\ : LocalMux
    port map (
            O => \N__39625\,
            I => \N__39611\
        );

    \I__8678\ : Span12Mux_s11_h
    port map (
            O => \N__39622\,
            I => \N__39611\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__39619\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8676\ : Odrv12
    port map (
            O => \N__39616\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8675\ : Odrv12
    port map (
            O => \N__39611\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__39604\,
            I => \N__39601\
        );

    \I__8673\ : InMux
    port map (
            O => \N__39601\,
            I => \N__39598\
        );

    \I__8672\ : LocalMux
    port map (
            O => \N__39598\,
            I => \N__39594\
        );

    \I__8671\ : InMux
    port map (
            O => \N__39597\,
            I => \N__39591\
        );

    \I__8670\ : Span4Mux_h
    port map (
            O => \N__39594\,
            I => \N__39588\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__39591\,
            I => \N__39585\
        );

    \I__8668\ : Span4Mux_h
    port map (
            O => \N__39588\,
            I => \N__39580\
        );

    \I__8667\ : Span4Mux_h
    port map (
            O => \N__39585\,
            I => \N__39576\
        );

    \I__8666\ : InMux
    port map (
            O => \N__39584\,
            I => \N__39573\
        );

    \I__8665\ : InMux
    port map (
            O => \N__39583\,
            I => \N__39570\
        );

    \I__8664\ : Span4Mux_v
    port map (
            O => \N__39580\,
            I => \N__39567\
        );

    \I__8663\ : InMux
    port map (
            O => \N__39579\,
            I => \N__39564\
        );

    \I__8662\ : Odrv4
    port map (
            O => \N__39576\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__39573\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__39570\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8659\ : Odrv4
    port map (
            O => \N__39567\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__39564\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__8657\ : InMux
    port map (
            O => \N__39553\,
            I => \N__39550\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__39550\,
            I => \N__39546\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39549\,
            I => \N__39542\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__39546\,
            I => \N__39539\
        );

    \I__8653\ : InMux
    port map (
            O => \N__39545\,
            I => \N__39536\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__39542\,
            I => \N__39533\
        );

    \I__8651\ : Span4Mux_h
    port map (
            O => \N__39539\,
            I => \N__39530\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__39536\,
            I => \N__39525\
        );

    \I__8649\ : Span4Mux_v
    port map (
            O => \N__39533\,
            I => \N__39525\
        );

    \I__8648\ : Odrv4
    port map (
            O => \N__39530\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8647\ : Odrv4
    port map (
            O => \N__39525\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__8646\ : CEMux
    port map (
            O => \N__39520\,
            I => \N__39517\
        );

    \I__8645\ : LocalMux
    port map (
            O => \N__39517\,
            I => \N__39514\
        );

    \I__8644\ : Span4Mux_v
    port map (
            O => \N__39514\,
            I => \N__39511\
        );

    \I__8643\ : Span4Mux_h
    port map (
            O => \N__39511\,
            I => \N__39508\
        );

    \I__8642\ : Odrv4
    port map (
            O => \N__39508\,
            I => \phase_controller_inst1.N_221_0\
        );

    \I__8641\ : CascadeMux
    port map (
            O => \N__39505\,
            I => \delay_measurement_inst.delay_tr_timer.N_424_cascade_\
        );

    \I__8640\ : InMux
    port map (
            O => \N__39502\,
            I => \N__39499\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__39499\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\
        );

    \I__8638\ : InMux
    port map (
            O => \N__39496\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39493\,
            I => \N__39490\
        );

    \I__8636\ : LocalMux
    port map (
            O => \N__39490\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\
        );

    \I__8635\ : InMux
    port map (
            O => \N__39487\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__8634\ : InMux
    port map (
            O => \N__39484\,
            I => \N__39481\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__39481\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\
        );

    \I__8632\ : InMux
    port map (
            O => \N__39478\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__8631\ : InMux
    port map (
            O => \N__39475\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__8630\ : InMux
    port map (
            O => \N__39472\,
            I => \N__39469\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__39469\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\
        );

    \I__8628\ : InMux
    port map (
            O => \N__39466\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__8627\ : InMux
    port map (
            O => \N__39463\,
            I => \N__39460\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39460\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\
        );

    \I__8625\ : InMux
    port map (
            O => \N__39457\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__8624\ : InMux
    port map (
            O => \N__39454\,
            I => \N__39451\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__39451\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\
        );

    \I__8622\ : InMux
    port map (
            O => \N__39448\,
            I => \bfn_16_18_0_\
        );

    \I__8621\ : InMux
    port map (
            O => \N__39445\,
            I => \N__39442\
        );

    \I__8620\ : LocalMux
    port map (
            O => \N__39442\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\
        );

    \I__8619\ : InMux
    port map (
            O => \N__39439\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__8618\ : InMux
    port map (
            O => \N__39436\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__8617\ : InMux
    port map (
            O => \N__39433\,
            I => \N__39430\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__39430\,
            I => \N__39427\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__39427\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\
        );

    \I__8614\ : InMux
    port map (
            O => \N__39424\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__8613\ : InMux
    port map (
            O => \N__39421\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__8612\ : InMux
    port map (
            O => \N__39418\,
            I => \N__39415\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__39415\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\
        );

    \I__8610\ : InMux
    port map (
            O => \N__39412\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__8609\ : InMux
    port map (
            O => \N__39409\,
            I => \N__39406\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__39406\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\
        );

    \I__8607\ : InMux
    port map (
            O => \N__39403\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__8606\ : InMux
    port map (
            O => \N__39400\,
            I => \N__39397\
        );

    \I__8605\ : LocalMux
    port map (
            O => \N__39397\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\
        );

    \I__8604\ : InMux
    port map (
            O => \N__39394\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__8603\ : InMux
    port map (
            O => \N__39391\,
            I => \N__39388\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__39388\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\
        );

    \I__8601\ : InMux
    port map (
            O => \N__39385\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__8600\ : InMux
    port map (
            O => \N__39382\,
            I => \N__39379\
        );

    \I__8599\ : LocalMux
    port map (
            O => \N__39379\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\
        );

    \I__8598\ : InMux
    port map (
            O => \N__39376\,
            I => \bfn_16_17_0_\
        );

    \I__8597\ : InMux
    port map (
            O => \N__39373\,
            I => \N__39370\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__39370\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\
        );

    \I__8595\ : InMux
    port map (
            O => \N__39367\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__8594\ : InMux
    port map (
            O => \N__39364\,
            I => \N__39361\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__39361\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39358\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__8591\ : InMux
    port map (
            O => \N__39355\,
            I => \N__39352\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__39352\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\
        );

    \I__8589\ : InMux
    port map (
            O => \N__39349\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__8588\ : InMux
    port map (
            O => \N__39346\,
            I => \N__39343\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__39343\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\
        );

    \I__8586\ : InMux
    port map (
            O => \N__39340\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__8585\ : InMux
    port map (
            O => \N__39337\,
            I => \N__39334\
        );

    \I__8584\ : LocalMux
    port map (
            O => \N__39334\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\
        );

    \I__8583\ : InMux
    port map (
            O => \N__39331\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__8582\ : InMux
    port map (
            O => \N__39328\,
            I => \N__39325\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__39325\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\
        );

    \I__8580\ : InMux
    port map (
            O => \N__39322\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__8579\ : InMux
    port map (
            O => \N__39319\,
            I => \N__39316\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__39316\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\
        );

    \I__8577\ : InMux
    port map (
            O => \N__39313\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__8576\ : InMux
    port map (
            O => \N__39310\,
            I => \N__39307\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39307\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\
        );

    \I__8574\ : InMux
    port map (
            O => \N__39304\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39301\,
            I => \N__39298\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__39298\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\
        );

    \I__8571\ : InMux
    port map (
            O => \N__39295\,
            I => \bfn_16_16_0_\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39292\,
            I => \N__39289\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__39289\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\
        );

    \I__8568\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39283\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__39283\,
            I => \N__39280\
        );

    \I__8566\ : Span4Mux_v
    port map (
            O => \N__39280\,
            I => \N__39276\
        );

    \I__8565\ : InMux
    port map (
            O => \N__39279\,
            I => \N__39273\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__39276\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__39273\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__39268\,
            I => \N__39265\
        );

    \I__8561\ : InMux
    port map (
            O => \N__39265\,
            I => \N__39262\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39262\,
            I => \N__39258\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__39261\,
            I => \N__39255\
        );

    \I__8558\ : Span4Mux_h
    port map (
            O => \N__39258\,
            I => \N__39252\
        );

    \I__8557\ : InMux
    port map (
            O => \N__39255\,
            I => \N__39249\
        );

    \I__8556\ : Odrv4
    port map (
            O => \N__39252\,
            I => measured_delay_tr_1
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39249\,
            I => measured_delay_tr_1
        );

    \I__8554\ : CascadeMux
    port map (
            O => \N__39244\,
            I => \N__39241\
        );

    \I__8553\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39238\
        );

    \I__8552\ : LocalMux
    port map (
            O => \N__39238\,
            I => \N__39235\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__39235\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__39232\,
            I => \N__39229\
        );

    \I__8549\ : InMux
    port map (
            O => \N__39229\,
            I => \N__39226\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__39226\,
            I => \N__39223\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__39223\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__8546\ : CascadeMux
    port map (
            O => \N__39220\,
            I => \N__39216\
        );

    \I__8545\ : CascadeMux
    port map (
            O => \N__39219\,
            I => \N__39211\
        );

    \I__8544\ : InMux
    port map (
            O => \N__39216\,
            I => \N__39208\
        );

    \I__8543\ : InMux
    port map (
            O => \N__39215\,
            I => \N__39205\
        );

    \I__8542\ : InMux
    port map (
            O => \N__39214\,
            I => \N__39200\
        );

    \I__8541\ : InMux
    port map (
            O => \N__39211\,
            I => \N__39200\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__39208\,
            I => \N__39197\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__39205\,
            I => \N__39192\
        );

    \I__8538\ : LocalMux
    port map (
            O => \N__39200\,
            I => \N__39192\
        );

    \I__8537\ : Span4Mux_v
    port map (
            O => \N__39197\,
            I => \N__39189\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__39192\,
            I => \N__39186\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__39189\,
            I => measured_delay_tr_9
        );

    \I__8534\ : Odrv4
    port map (
            O => \N__39186\,
            I => measured_delay_tr_9
        );

    \I__8533\ : InMux
    port map (
            O => \N__39181\,
            I => \N__39178\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__39178\,
            I => \N__39175\
        );

    \I__8531\ : Span4Mux_v
    port map (
            O => \N__39175\,
            I => \N__39172\
        );

    \I__8530\ : Span4Mux_h
    port map (
            O => \N__39172\,
            I => \N__39169\
        );

    \I__8529\ : Odrv4
    port map (
            O => \N__39169\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3\
        );

    \I__8528\ : InMux
    port map (
            O => \N__39166\,
            I => \N__39161\
        );

    \I__8527\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39156\
        );

    \I__8526\ : InMux
    port map (
            O => \N__39164\,
            I => \N__39156\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__39161\,
            I => \N__39151\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__39156\,
            I => \N__39151\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__39151\,
            I => \N__39147\
        );

    \I__8522\ : CascadeMux
    port map (
            O => \N__39150\,
            I => \N__39143\
        );

    \I__8521\ : Span4Mux_h
    port map (
            O => \N__39147\,
            I => \N__39140\
        );

    \I__8520\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39135\
        );

    \I__8519\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39135\
        );

    \I__8518\ : Odrv4
    port map (
            O => \N__39140\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__39135\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\
        );

    \I__8516\ : InMux
    port map (
            O => \N__39130\,
            I => \N__39124\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39129\,
            I => \N__39124\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__39124\,
            I => \N__39119\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39123\,
            I => \N__39116\
        );

    \I__8512\ : CascadeMux
    port map (
            O => \N__39122\,
            I => \N__39113\
        );

    \I__8511\ : Span4Mux_v
    port map (
            O => \N__39119\,
            I => \N__39107\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__39116\,
            I => \N__39107\
        );

    \I__8509\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39102\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39102\
        );

    \I__8507\ : Span4Mux_h
    port map (
            O => \N__39107\,
            I => \N__39099\
        );

    \I__8506\ : LocalMux
    port map (
            O => \N__39102\,
            I => measured_delay_tr_3
        );

    \I__8505\ : Odrv4
    port map (
            O => \N__39099\,
            I => measured_delay_tr_3
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__39094\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_\
        );

    \I__8503\ : InMux
    port map (
            O => \N__39091\,
            I => \N__39082\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39082\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39082\
        );

    \I__8500\ : LocalMux
    port map (
            O => \N__39082\,
            I => \N__39076\
        );

    \I__8499\ : InMux
    port map (
            O => \N__39081\,
            I => \N__39069\
        );

    \I__8498\ : InMux
    port map (
            O => \N__39080\,
            I => \N__39069\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39079\,
            I => \N__39069\
        );

    \I__8496\ : Span12Mux_h
    port map (
            O => \N__39076\,
            I => \N__39066\
        );

    \I__8495\ : LocalMux
    port map (
            O => \N__39069\,
            I => \N__39063\
        );

    \I__8494\ : Odrv12
    port map (
            O => \N__39066\,
            I => \phase_controller_inst1.stoper_tr.N_20_li\
        );

    \I__8493\ : Odrv12
    port map (
            O => \N__39063\,
            I => \phase_controller_inst1.stoper_tr.N_20_li\
        );

    \I__8492\ : CascadeMux
    port map (
            O => \N__39058\,
            I => \N__39055\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39055\,
            I => \N__39052\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__39052\,
            I => \N__39049\
        );

    \I__8489\ : Odrv12
    port map (
            O => \N__39049\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__8488\ : InMux
    port map (
            O => \N__39046\,
            I => \N__39042\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39045\,
            I => \N__39039\
        );

    \I__8486\ : LocalMux
    port map (
            O => \N__39042\,
            I => \N__39034\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39039\,
            I => \N__39031\
        );

    \I__8484\ : CascadeMux
    port map (
            O => \N__39038\,
            I => \N__39028\
        );

    \I__8483\ : InMux
    port map (
            O => \N__39037\,
            I => \N__39025\
        );

    \I__8482\ : Span4Mux_v
    port map (
            O => \N__39034\,
            I => \N__39022\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__39031\,
            I => \N__39019\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39028\,
            I => \N__39016\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__39025\,
            I => \N__39011\
        );

    \I__8478\ : Span4Mux_h
    port map (
            O => \N__39022\,
            I => \N__39011\
        );

    \I__8477\ : Odrv4
    port map (
            O => \N__39019\,
            I => measured_delay_tr_8
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39016\,
            I => measured_delay_tr_8
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__39011\,
            I => measured_delay_tr_8
        );

    \I__8474\ : InMux
    port map (
            O => \N__39004\,
            I => \N__38999\
        );

    \I__8473\ : InMux
    port map (
            O => \N__39003\,
            I => \N__38995\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39002\,
            I => \N__38992\
        );

    \I__8471\ : LocalMux
    port map (
            O => \N__38999\,
            I => \N__38989\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__38998\,
            I => \N__38986\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__38995\,
            I => \N__38983\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__38992\,
            I => \N__38980\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__38989\,
            I => \N__38977\
        );

    \I__8466\ : InMux
    port map (
            O => \N__38986\,
            I => \N__38974\
        );

    \I__8465\ : Span4Mux_v
    port map (
            O => \N__38983\,
            I => \N__38969\
        );

    \I__8464\ : Span4Mux_h
    port map (
            O => \N__38980\,
            I => \N__38969\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__38977\,
            I => measured_delay_tr_7
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__38974\,
            I => measured_delay_tr_7
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__38969\,
            I => measured_delay_tr_7
        );

    \I__8460\ : InMux
    port map (
            O => \N__38962\,
            I => \N__38959\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__38959\,
            I => \N__38956\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__38956\,
            I => \N__38951\
        );

    \I__8457\ : InMux
    port map (
            O => \N__38955\,
            I => \N__38948\
        );

    \I__8456\ : InMux
    port map (
            O => \N__38954\,
            I => \N__38945\
        );

    \I__8455\ : Span4Mux_h
    port map (
            O => \N__38951\,
            I => \N__38942\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__38948\,
            I => \N__38937\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__38945\,
            I => \N__38937\
        );

    \I__8452\ : Sp12to4
    port map (
            O => \N__38942\,
            I => \N__38934\
        );

    \I__8451\ : Span4Mux_v
    port map (
            O => \N__38937\,
            I => \N__38931\
        );

    \I__8450\ : Odrv12
    port map (
            O => \N__38934\,
            I => measured_delay_tr_6
        );

    \I__8449\ : Odrv4
    port map (
            O => \N__38931\,
            I => measured_delay_tr_6
        );

    \I__8448\ : CascadeMux
    port map (
            O => \N__38926\,
            I => \N__38923\
        );

    \I__8447\ : InMux
    port map (
            O => \N__38923\,
            I => \N__38920\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__38920\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\
        );

    \I__8445\ : CascadeMux
    port map (
            O => \N__38917\,
            I => \N__38914\
        );

    \I__8444\ : InMux
    port map (
            O => \N__38914\,
            I => \N__38909\
        );

    \I__8443\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38906\
        );

    \I__8442\ : CascadeMux
    port map (
            O => \N__38912\,
            I => \N__38903\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__38909\,
            I => \N__38898\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__38906\,
            I => \N__38898\
        );

    \I__8439\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38893\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__38898\,
            I => \N__38890\
        );

    \I__8437\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38885\
        );

    \I__8436\ : InMux
    port map (
            O => \N__38896\,
            I => \N__38885\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__38893\,
            I => \N__38876\
        );

    \I__8434\ : Span4Mux_h
    port map (
            O => \N__38890\,
            I => \N__38876\
        );

    \I__8433\ : LocalMux
    port map (
            O => \N__38885\,
            I => \N__38876\
        );

    \I__8432\ : InMux
    port map (
            O => \N__38884\,
            I => \N__38873\
        );

    \I__8431\ : CascadeMux
    port map (
            O => \N__38883\,
            I => \N__38870\
        );

    \I__8430\ : Span4Mux_h
    port map (
            O => \N__38876\,
            I => \N__38864\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__38873\,
            I => \N__38861\
        );

    \I__8428\ : InMux
    port map (
            O => \N__38870\,
            I => \N__38858\
        );

    \I__8427\ : InMux
    port map (
            O => \N__38869\,
            I => \N__38851\
        );

    \I__8426\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38851\
        );

    \I__8425\ : InMux
    port map (
            O => \N__38867\,
            I => \N__38851\
        );

    \I__8424\ : Span4Mux_v
    port map (
            O => \N__38864\,
            I => \N__38848\
        );

    \I__8423\ : Span4Mux_h
    port map (
            O => \N__38861\,
            I => \N__38845\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__38858\,
            I => measured_delay_tr_15
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__38851\,
            I => measured_delay_tr_15
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__38848\,
            I => measured_delay_tr_15
        );

    \I__8419\ : Odrv4
    port map (
            O => \N__38845\,
            I => measured_delay_tr_15
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__38836\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_\
        );

    \I__8417\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38830\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__38830\,
            I => \N__38827\
        );

    \I__8415\ : Span4Mux_h
    port map (
            O => \N__38827\,
            I => \N__38820\
        );

    \I__8414\ : InMux
    port map (
            O => \N__38826\,
            I => \N__38815\
        );

    \I__8413\ : InMux
    port map (
            O => \N__38825\,
            I => \N__38815\
        );

    \I__8412\ : InMux
    port map (
            O => \N__38824\,
            I => \N__38810\
        );

    \I__8411\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38810\
        );

    \I__8410\ : Span4Mux_v
    port map (
            O => \N__38820\,
            I => \N__38805\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__38815\,
            I => \N__38805\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__38810\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__38805\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\
        );

    \I__8406\ : InMux
    port map (
            O => \N__38800\,
            I => \N__38795\
        );

    \I__8405\ : CascadeMux
    port map (
            O => \N__38799\,
            I => \N__38792\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__38798\,
            I => \N__38789\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38795\,
            I => \N__38786\
        );

    \I__8402\ : InMux
    port map (
            O => \N__38792\,
            I => \N__38783\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38780\
        );

    \I__8400\ : Span4Mux_v
    port map (
            O => \N__38786\,
            I => \N__38777\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__38783\,
            I => \N__38772\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38780\,
            I => \N__38772\
        );

    \I__8397\ : Span4Mux_h
    port map (
            O => \N__38777\,
            I => \N__38769\
        );

    \I__8396\ : Span4Mux_h
    port map (
            O => \N__38772\,
            I => \N__38766\
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__38769\,
            I => measured_delay_tr_5
        );

    \I__8394\ : Odrv4
    port map (
            O => \N__38766\,
            I => measured_delay_tr_5
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__38761\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__38758\,
            I => \N__38755\
        );

    \I__8391\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38752\
        );

    \I__8390\ : LocalMux
    port map (
            O => \N__38752\,
            I => \N__38749\
        );

    \I__8389\ : Span4Mux_h
    port map (
            O => \N__38749\,
            I => \N__38746\
        );

    \I__8388\ : Odrv4
    port map (
            O => \N__38746\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__8387\ : InMux
    port map (
            O => \N__38743\,
            I => \N__38740\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__38740\,
            I => \N__38737\
        );

    \I__8385\ : Odrv12
    port map (
            O => \N__38737\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\
        );

    \I__8384\ : InMux
    port map (
            O => \N__38734\,
            I => \N__38730\
        );

    \I__8383\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38727\
        );

    \I__8382\ : LocalMux
    port map (
            O => \N__38730\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8381\ : LocalMux
    port map (
            O => \N__38727\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8380\ : CascadeMux
    port map (
            O => \N__38722\,
            I => \N__38719\
        );

    \I__8379\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38716\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__38716\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38709\
        );

    \I__8376\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38706\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__38709\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__38706\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8373\ : InMux
    port map (
            O => \N__38701\,
            I => \N__38698\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__38698\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__38695\,
            I => \N__38692\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38688\
        );

    \I__8369\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38685\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__38688\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__38685\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38680\,
            I => \N__38677\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__38677\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__8364\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38670\
        );

    \I__8363\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38667\
        );

    \I__8362\ : LocalMux
    port map (
            O => \N__38670\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__38667\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38662\,
            I => \N__38659\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__38659\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__8358\ : InMux
    port map (
            O => \N__38656\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8357\ : CascadeMux
    port map (
            O => \N__38653\,
            I => \N__38650\
        );

    \I__8356\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38647\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__38647\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__38644\,
            I => \N__38641\
        );

    \I__8353\ : InMux
    port map (
            O => \N__38641\,
            I => \N__38638\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38638\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__8351\ : CascadeMux
    port map (
            O => \N__38635\,
            I => \N__38632\
        );

    \I__8350\ : InMux
    port map (
            O => \N__38632\,
            I => \N__38629\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__38629\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__8348\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38623\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__38623\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__8346\ : CascadeMux
    port map (
            O => \N__38620\,
            I => \N__38617\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38617\,
            I => \N__38614\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__38614\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__8343\ : InMux
    port map (
            O => \N__38611\,
            I => \N__38607\
        );

    \I__8342\ : InMux
    port map (
            O => \N__38610\,
            I => \N__38604\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__38607\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__38604\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8339\ : InMux
    port map (
            O => \N__38599\,
            I => \N__38596\
        );

    \I__8338\ : LocalMux
    port map (
            O => \N__38596\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__8337\ : CascadeMux
    port map (
            O => \N__38593\,
            I => \N__38590\
        );

    \I__8336\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38587\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__38587\,
            I => \N__38584\
        );

    \I__8334\ : Odrv4
    port map (
            O => \N__38584\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__38581\,
            I => \N__38578\
        );

    \I__8332\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38574\
        );

    \I__8331\ : InMux
    port map (
            O => \N__38577\,
            I => \N__38571\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__38574\,
            I => \N__38568\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38565\
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__38568\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8327\ : Odrv4
    port map (
            O => \N__38565\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8326\ : InMux
    port map (
            O => \N__38560\,
            I => \N__38557\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__38557\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__8324\ : CascadeMux
    port map (
            O => \N__38554\,
            I => \N__38551\
        );

    \I__8323\ : InMux
    port map (
            O => \N__38551\,
            I => \N__38548\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__38548\,
            I => \N__38545\
        );

    \I__8321\ : Odrv4
    port map (
            O => \N__38545\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__8320\ : InMux
    port map (
            O => \N__38542\,
            I => \N__38539\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__38539\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__8318\ : CascadeMux
    port map (
            O => \N__38536\,
            I => \N__38533\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38533\,
            I => \N__38530\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__38530\,
            I => \N__38527\
        );

    \I__8315\ : Odrv4
    port map (
            O => \N__38527\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__8314\ : InMux
    port map (
            O => \N__38524\,
            I => \N__38520\
        );

    \I__8313\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38517\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__38520\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8311\ : LocalMux
    port map (
            O => \N__38517\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8310\ : InMux
    port map (
            O => \N__38512\,
            I => \N__38509\
        );

    \I__8309\ : LocalMux
    port map (
            O => \N__38509\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__8308\ : CascadeMux
    port map (
            O => \N__38506\,
            I => \N__38503\
        );

    \I__8307\ : InMux
    port map (
            O => \N__38503\,
            I => \N__38499\
        );

    \I__8306\ : InMux
    port map (
            O => \N__38502\,
            I => \N__38496\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__38499\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__38496\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8303\ : CascadeMux
    port map (
            O => \N__38491\,
            I => \N__38488\
        );

    \I__8302\ : InMux
    port map (
            O => \N__38488\,
            I => \N__38485\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__38485\,
            I => \N__38482\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__38482\,
            I => \N__38479\
        );

    \I__8299\ : Odrv4
    port map (
            O => \N__38479\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__8298\ : InMux
    port map (
            O => \N__38476\,
            I => \N__38473\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__38473\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__8296\ : CascadeMux
    port map (
            O => \N__38470\,
            I => \N__38467\
        );

    \I__8295\ : InMux
    port map (
            O => \N__38467\,
            I => \N__38464\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__38464\,
            I => \N__38461\
        );

    \I__8293\ : Odrv4
    port map (
            O => \N__38461\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38454\
        );

    \I__8291\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38451\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__38454\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__38451\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38446\,
            I => \N__38443\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__38443\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__38440\,
            I => \N__38437\
        );

    \I__8285\ : InMux
    port map (
            O => \N__38437\,
            I => \N__38434\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38434\,
            I => \N__38431\
        );

    \I__8283\ : Span4Mux_v
    port map (
            O => \N__38431\,
            I => \N__38428\
        );

    \I__8282\ : Odrv4
    port map (
            O => \N__38428\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__8281\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38421\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38424\,
            I => \N__38418\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38421\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__38418\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8277\ : InMux
    port map (
            O => \N__38413\,
            I => \N__38410\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__38410\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__38407\,
            I => \N__38403\
        );

    \I__8274\ : InMux
    port map (
            O => \N__38406\,
            I => \N__38399\
        );

    \I__8273\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38396\
        );

    \I__8272\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38393\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__38399\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38396\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__38393\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8268\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38383\
        );

    \I__8267\ : LocalMux
    port map (
            O => \N__38383\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38380\,
            I => \N__38376\
        );

    \I__8265\ : InMux
    port map (
            O => \N__38379\,
            I => \N__38373\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__38376\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38373\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8262\ : InMux
    port map (
            O => \N__38368\,
            I => \N__38365\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__38365\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__38362\,
            I => \N__38359\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38355\
        );

    \I__8258\ : InMux
    port map (
            O => \N__38358\,
            I => \N__38352\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__38355\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__38352\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8255\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38344\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__38344\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__8253\ : CascadeMux
    port map (
            O => \N__38341\,
            I => \N__38338\
        );

    \I__8252\ : InMux
    port map (
            O => \N__38338\,
            I => \N__38335\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__38335\,
            I => \N__38332\
        );

    \I__8250\ : Odrv4
    port map (
            O => \N__38332\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__8249\ : InMux
    port map (
            O => \N__38329\,
            I => \N__38325\
        );

    \I__8248\ : InMux
    port map (
            O => \N__38328\,
            I => \N__38322\
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__38325\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__38322\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38314\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38314\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__8243\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38307\
        );

    \I__8242\ : InMux
    port map (
            O => \N__38310\,
            I => \N__38304\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__38307\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__38304\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8239\ : InMux
    port map (
            O => \N__38299\,
            I => \N__38296\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__38296\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__8237\ : CascadeMux
    port map (
            O => \N__38293\,
            I => \N__38290\
        );

    \I__8236\ : InMux
    port map (
            O => \N__38290\,
            I => \N__38287\
        );

    \I__8235\ : LocalMux
    port map (
            O => \N__38287\,
            I => \N__38284\
        );

    \I__8234\ : Odrv4
    port map (
            O => \N__38284\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\
        );

    \I__8233\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38277\
        );

    \I__8232\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38274\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38277\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__38274\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38269\,
            I => \N__38266\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38266\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__8227\ : CascadeMux
    port map (
            O => \N__38263\,
            I => \N__38260\
        );

    \I__8226\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38257\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38254\
        );

    \I__8224\ : Odrv4
    port map (
            O => \N__38254\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__8223\ : InMux
    port map (
            O => \N__38251\,
            I => \N__38247\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38250\,
            I => \N__38244\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__38247\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__38244\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38239\,
            I => \N__38236\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__38236\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__38233\,
            I => \N__38230\
        );

    \I__8216\ : InMux
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__8215\ : LocalMux
    port map (
            O => \N__38227\,
            I => \N__38224\
        );

    \I__8214\ : Span4Mux_h
    port map (
            O => \N__38224\,
            I => \N__38221\
        );

    \I__8213\ : Odrv4
    port map (
            O => \N__38221\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__8212\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38214\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38211\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__38214\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__38211\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__38206\,
            I => \N__38203\
        );

    \I__8207\ : InMux
    port map (
            O => \N__38203\,
            I => \N__38200\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__38200\,
            I => \N__38197\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__38197\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38194\,
            I => \N__38191\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38191\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__38188\,
            I => \N__38185\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38185\,
            I => \N__38182\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__38182\,
            I => \N__38179\
        );

    \I__8199\ : Odrv12
    port map (
            O => \N__38179\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38176\,
            I => \N__38173\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38173\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__8196\ : CascadeMux
    port map (
            O => \N__38170\,
            I => \N__38167\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38167\,
            I => \N__38164\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38164\,
            I => \N__38161\
        );

    \I__8193\ : Odrv4
    port map (
            O => \N__38161\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__8192\ : InMux
    port map (
            O => \N__38158\,
            I => \N__38155\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__38155\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__38152\,
            I => \N__38149\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38149\,
            I => \N__38146\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__38146\,
            I => \N__38143\
        );

    \I__8187\ : Odrv4
    port map (
            O => \N__38143\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38140\,
            I => \N__38137\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38137\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__8184\ : CascadeMux
    port map (
            O => \N__38134\,
            I => \N__38131\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38128\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__38128\,
            I => \N__38125\
        );

    \I__8181\ : Span4Mux_h
    port map (
            O => \N__38125\,
            I => \N__38122\
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__38122\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__38116\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38113\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__8176\ : CascadeMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38107\,
            I => \N__38104\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38101\
        );

    \I__8173\ : Odrv4
    port map (
            O => \N__38101\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__8172\ : InMux
    port map (
            O => \N__38098\,
            I => \N__38095\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38095\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__8170\ : CascadeMux
    port map (
            O => \N__38092\,
            I => \N__38089\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38089\,
            I => \N__38086\
        );

    \I__8168\ : LocalMux
    port map (
            O => \N__38086\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38080\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38080\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__8165\ : CascadeMux
    port map (
            O => \N__38077\,
            I => \N__38074\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38074\,
            I => \N__38071\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__38071\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38068\,
            I => \N__38065\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38065\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__38062\,
            I => \N__38059\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38059\,
            I => \N__38056\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38056\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__8157\ : InMux
    port map (
            O => \N__38053\,
            I => \N__38050\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__38050\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__38047\,
            I => \N__38044\
        );

    \I__8154\ : InMux
    port map (
            O => \N__38044\,
            I => \N__38041\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38041\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38035\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__38035\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__38032\,
            I => \N__38029\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38029\,
            I => \N__38026\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__38026\,
            I => \N__38023\
        );

    \I__8147\ : Odrv12
    port map (
            O => \N__38023\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38020\,
            I => \N__38017\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__38017\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__8144\ : CascadeMux
    port map (
            O => \N__38014\,
            I => \N__38011\
        );

    \I__8143\ : InMux
    port map (
            O => \N__38011\,
            I => \N__38008\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__38008\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38005\,
            I => \N__38002\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__38002\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__8139\ : CascadeMux
    port map (
            O => \N__37999\,
            I => \N__37996\
        );

    \I__8138\ : InMux
    port map (
            O => \N__37996\,
            I => \N__37993\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__37993\,
            I => \N__37990\
        );

    \I__8136\ : Span4Mux_v
    port map (
            O => \N__37990\,
            I => \N__37987\
        );

    \I__8135\ : Span4Mux_h
    port map (
            O => \N__37987\,
            I => \N__37984\
        );

    \I__8134\ : Odrv4
    port map (
            O => \N__37984\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__8133\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37978\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__37978\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__8131\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37972\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__37972\,
            I => \N__37969\
        );

    \I__8129\ : Odrv4
    port map (
            O => \N__37969\,
            I => delay_hc_input_c
        );

    \I__8128\ : InMux
    port map (
            O => \N__37966\,
            I => \N__37963\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__37963\,
            I => \N__37960\
        );

    \I__8126\ : Odrv12
    port map (
            O => \N__37960\,
            I => delay_hc_d1
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__37957\,
            I => \N__37954\
        );

    \I__8124\ : InMux
    port map (
            O => \N__37954\,
            I => \N__37951\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__37951\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\
        );

    \I__8122\ : InMux
    port map (
            O => \N__37948\,
            I => \N__37945\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__37945\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__8120\ : CascadeMux
    port map (
            O => \N__37942\,
            I => \N__37939\
        );

    \I__8119\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37936\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__37936\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__8117\ : CascadeMux
    port map (
            O => \N__37933\,
            I => \N__37930\
        );

    \I__8116\ : InMux
    port map (
            O => \N__37930\,
            I => \N__37927\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__37927\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__8114\ : InMux
    port map (
            O => \N__37924\,
            I => \N__37921\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__37921\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__8112\ : CascadeMux
    port map (
            O => \N__37918\,
            I => \N__37915\
        );

    \I__8111\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37912\
        );

    \I__8110\ : LocalMux
    port map (
            O => \N__37912\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__8109\ : InMux
    port map (
            O => \N__37909\,
            I => \N__37906\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__37906\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__8107\ : CascadeMux
    port map (
            O => \N__37903\,
            I => \N__37900\
        );

    \I__8106\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37897\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__37897\,
            I => \N__37894\
        );

    \I__8104\ : Odrv4
    port map (
            O => \N__37894\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__8103\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37888\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__37888\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__8101\ : CascadeMux
    port map (
            O => \N__37885\,
            I => \N__37882\
        );

    \I__8100\ : InMux
    port map (
            O => \N__37882\,
            I => \N__37879\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__37879\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__8098\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37873\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__37873\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__8096\ : CascadeMux
    port map (
            O => \N__37870\,
            I => \N__37867\
        );

    \I__8095\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37864\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__37864\,
            I => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\
        );

    \I__8093\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37858\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__37858\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__8091\ : CascadeMux
    port map (
            O => \N__37855\,
            I => \N__37852\
        );

    \I__8090\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37849\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__37849\,
            I => \N__37846\
        );

    \I__8088\ : Span4Mux_v
    port map (
            O => \N__37846\,
            I => \N__37843\
        );

    \I__8087\ : Odrv4
    port map (
            O => \N__37843\,
            I => \current_shift_inst.z_5_23\
        );

    \I__8086\ : InMux
    port map (
            O => \N__37840\,
            I => \current_shift_inst.z_5_cry_22\
        );

    \I__8085\ : CascadeMux
    port map (
            O => \N__37837\,
            I => \N__37834\
        );

    \I__8084\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37831\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__37831\,
            I => \N__37828\
        );

    \I__8082\ : Span4Mux_h
    port map (
            O => \N__37828\,
            I => \N__37825\
        );

    \I__8081\ : Odrv4
    port map (
            O => \N__37825\,
            I => \current_shift_inst.z_5_24\
        );

    \I__8080\ : InMux
    port map (
            O => \N__37822\,
            I => \current_shift_inst.z_5_cry_23\
        );

    \I__8079\ : InMux
    port map (
            O => \N__37819\,
            I => \N__37816\
        );

    \I__8078\ : LocalMux
    port map (
            O => \N__37816\,
            I => \N__37813\
        );

    \I__8077\ : Span4Mux_v
    port map (
            O => \N__37813\,
            I => \N__37810\
        );

    \I__8076\ : Odrv4
    port map (
            O => \N__37810\,
            I => \current_shift_inst.z_5_25\
        );

    \I__8075\ : InMux
    port map (
            O => \N__37807\,
            I => \bfn_15_24_0_\
        );

    \I__8074\ : CascadeMux
    port map (
            O => \N__37804\,
            I => \N__37801\
        );

    \I__8073\ : InMux
    port map (
            O => \N__37801\,
            I => \N__37798\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__37798\,
            I => \N__37795\
        );

    \I__8071\ : Span4Mux_h
    port map (
            O => \N__37795\,
            I => \N__37792\
        );

    \I__8070\ : Odrv4
    port map (
            O => \N__37792\,
            I => \current_shift_inst.z_5_26\
        );

    \I__8069\ : InMux
    port map (
            O => \N__37789\,
            I => \current_shift_inst.z_5_cry_25\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__37786\,
            I => \N__37783\
        );

    \I__8067\ : InMux
    port map (
            O => \N__37783\,
            I => \N__37780\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__37780\,
            I => \N__37777\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__37777\,
            I => \N__37774\
        );

    \I__8064\ : Odrv4
    port map (
            O => \N__37774\,
            I => \current_shift_inst.z_5_27\
        );

    \I__8063\ : InMux
    port map (
            O => \N__37771\,
            I => \current_shift_inst.z_5_cry_26\
        );

    \I__8062\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37765\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__37765\,
            I => \N__37762\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__37762\,
            I => \N__37759\
        );

    \I__8059\ : Odrv4
    port map (
            O => \N__37759\,
            I => \current_shift_inst.z_5_28\
        );

    \I__8058\ : InMux
    port map (
            O => \N__37756\,
            I => \current_shift_inst.z_5_cry_27\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__37753\,
            I => \N__37750\
        );

    \I__8056\ : InMux
    port map (
            O => \N__37750\,
            I => \N__37747\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__37747\,
            I => \N__37744\
        );

    \I__8054\ : Span4Mux_v
    port map (
            O => \N__37744\,
            I => \N__37741\
        );

    \I__8053\ : Odrv4
    port map (
            O => \N__37741\,
            I => \current_shift_inst.z_5_29\
        );

    \I__8052\ : InMux
    port map (
            O => \N__37738\,
            I => \current_shift_inst.z_5_cry_28\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37732\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__37732\,
            I => \N__37729\
        );

    \I__8049\ : Span4Mux_v
    port map (
            O => \N__37729\,
            I => \N__37726\
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__37726\,
            I => \current_shift_inst.z_5_30\
        );

    \I__8047\ : InMux
    port map (
            O => \N__37723\,
            I => \current_shift_inst.z_5_cry_29\
        );

    \I__8046\ : InMux
    port map (
            O => \N__37720\,
            I => \current_shift_inst.z_5_cry_30\
        );

    \I__8045\ : InMux
    port map (
            O => \N__37717\,
            I => \N__37714\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__37714\,
            I => \N__37711\
        );

    \I__8043\ : Span4Mux_v
    port map (
            O => \N__37711\,
            I => \N__37708\
        );

    \I__8042\ : Odrv4
    port map (
            O => \N__37708\,
            I => \current_shift_inst.z_5_cry_30_THRU_CO\
        );

    \I__8041\ : CascadeMux
    port map (
            O => \N__37705\,
            I => \N__37702\
        );

    \I__8040\ : InMux
    port map (
            O => \N__37702\,
            I => \N__37699\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37696\
        );

    \I__8038\ : Span4Mux_v
    port map (
            O => \N__37696\,
            I => \N__37693\
        );

    \I__8037\ : Odrv4
    port map (
            O => \N__37693\,
            I => \current_shift_inst.z_5_15\
        );

    \I__8036\ : InMux
    port map (
            O => \N__37690\,
            I => \current_shift_inst.z_5_cry_14\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__37687\,
            I => \N__37684\
        );

    \I__8034\ : InMux
    port map (
            O => \N__37684\,
            I => \N__37681\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__37681\,
            I => \N__37678\
        );

    \I__8032\ : Span4Mux_h
    port map (
            O => \N__37678\,
            I => \N__37675\
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__37675\,
            I => \current_shift_inst.z_5_16\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37672\,
            I => \current_shift_inst.z_5_cry_15\
        );

    \I__8029\ : InMux
    port map (
            O => \N__37669\,
            I => \N__37666\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__37666\,
            I => \N__37663\
        );

    \I__8027\ : Span4Mux_v
    port map (
            O => \N__37663\,
            I => \N__37660\
        );

    \I__8026\ : Odrv4
    port map (
            O => \N__37660\,
            I => \current_shift_inst.z_5_17\
        );

    \I__8025\ : InMux
    port map (
            O => \N__37657\,
            I => \bfn_15_23_0_\
        );

    \I__8024\ : CascadeMux
    port map (
            O => \N__37654\,
            I => \N__37651\
        );

    \I__8023\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37648\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__37648\,
            I => \N__37645\
        );

    \I__8021\ : Span4Mux_h
    port map (
            O => \N__37645\,
            I => \N__37642\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__37642\,
            I => \current_shift_inst.z_5_18\
        );

    \I__8019\ : InMux
    port map (
            O => \N__37639\,
            I => \current_shift_inst.z_5_cry_17\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37636\,
            I => \N__37633\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__37633\,
            I => \N__37630\
        );

    \I__8016\ : Odrv4
    port map (
            O => \N__37630\,
            I => \current_shift_inst.z_5_19\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37627\,
            I => \current_shift_inst.z_5_cry_18\
        );

    \I__8014\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37621\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__37621\,
            I => \N__37618\
        );

    \I__8012\ : Span4Mux_h
    port map (
            O => \N__37618\,
            I => \N__37615\
        );

    \I__8011\ : Odrv4
    port map (
            O => \N__37615\,
            I => \current_shift_inst.z_5_20\
        );

    \I__8010\ : InMux
    port map (
            O => \N__37612\,
            I => \current_shift_inst.z_5_cry_19\
        );

    \I__8009\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37606\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__37606\,
            I => \N__37603\
        );

    \I__8007\ : Odrv4
    port map (
            O => \N__37603\,
            I => \current_shift_inst.z_5_21\
        );

    \I__8006\ : InMux
    port map (
            O => \N__37600\,
            I => \current_shift_inst.z_5_cry_20\
        );

    \I__8005\ : InMux
    port map (
            O => \N__37597\,
            I => \N__37594\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__37594\,
            I => \N__37591\
        );

    \I__8003\ : Span4Mux_v
    port map (
            O => \N__37591\,
            I => \N__37588\
        );

    \I__8002\ : Odrv4
    port map (
            O => \N__37588\,
            I => \current_shift_inst.z_5_22\
        );

    \I__8001\ : InMux
    port map (
            O => \N__37585\,
            I => \current_shift_inst.z_5_cry_21\
        );

    \I__8000\ : CascadeMux
    port map (
            O => \N__37582\,
            I => \N__37579\
        );

    \I__7999\ : InMux
    port map (
            O => \N__37579\,
            I => \N__37576\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__37576\,
            I => \N__37573\
        );

    \I__7997\ : Span4Mux_v
    port map (
            O => \N__37573\,
            I => \N__37570\
        );

    \I__7996\ : Odrv4
    port map (
            O => \N__37570\,
            I => \current_shift_inst.z_5_7\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37567\,
            I => \current_shift_inst.z_5_cry_6\
        );

    \I__7994\ : InMux
    port map (
            O => \N__37564\,
            I => \N__37561\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__37561\,
            I => \N__37558\
        );

    \I__7992\ : Span4Mux_h
    port map (
            O => \N__37558\,
            I => \N__37555\
        );

    \I__7991\ : Odrv4
    port map (
            O => \N__37555\,
            I => \current_shift_inst.z_5_8\
        );

    \I__7990\ : InMux
    port map (
            O => \N__37552\,
            I => \current_shift_inst.z_5_cry_7\
        );

    \I__7989\ : CascadeMux
    port map (
            O => \N__37549\,
            I => \N__37546\
        );

    \I__7988\ : InMux
    port map (
            O => \N__37546\,
            I => \N__37543\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__37543\,
            I => \N__37540\
        );

    \I__7986\ : Odrv4
    port map (
            O => \N__37540\,
            I => \current_shift_inst.z_5_9\
        );

    \I__7985\ : InMux
    port map (
            O => \N__37537\,
            I => \bfn_15_22_0_\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37534\,
            I => \N__37531\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__37531\,
            I => \N__37528\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__37528\,
            I => \current_shift_inst.z_5_10\
        );

    \I__7981\ : InMux
    port map (
            O => \N__37525\,
            I => \current_shift_inst.z_5_cry_9\
        );

    \I__7980\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37519\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__37519\,
            I => \N__37516\
        );

    \I__7978\ : Odrv4
    port map (
            O => \N__37516\,
            I => \current_shift_inst.z_5_11\
        );

    \I__7977\ : InMux
    port map (
            O => \N__37513\,
            I => \current_shift_inst.z_5_cry_10\
        );

    \I__7976\ : CascadeMux
    port map (
            O => \N__37510\,
            I => \N__37507\
        );

    \I__7975\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37504\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__37504\,
            I => \N__37501\
        );

    \I__7973\ : Odrv4
    port map (
            O => \N__37501\,
            I => \current_shift_inst.z_5_12\
        );

    \I__7972\ : InMux
    port map (
            O => \N__37498\,
            I => \current_shift_inst.z_5_cry_11\
        );

    \I__7971\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37492\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__37492\,
            I => \N__37489\
        );

    \I__7969\ : Odrv4
    port map (
            O => \N__37489\,
            I => \current_shift_inst.z_5_13\
        );

    \I__7968\ : InMux
    port map (
            O => \N__37486\,
            I => \current_shift_inst.z_5_cry_12\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__37483\,
            I => \N__37480\
        );

    \I__7966\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37477\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__37477\,
            I => \N__37474\
        );

    \I__7964\ : Span4Mux_v
    port map (
            O => \N__37474\,
            I => \N__37471\
        );

    \I__7963\ : Odrv4
    port map (
            O => \N__37471\,
            I => \current_shift_inst.z_5_14\
        );

    \I__7962\ : InMux
    port map (
            O => \N__37468\,
            I => \current_shift_inst.z_5_cry_13\
        );

    \I__7961\ : InMux
    port map (
            O => \N__37465\,
            I => \N__37462\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__37462\,
            I => \N__37459\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__37459\,
            I => \N__37456\
        );

    \I__7958\ : Span4Mux_h
    port map (
            O => \N__37456\,
            I => \N__37453\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__37453\,
            I => \current_shift_inst.N_1742_i\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__37450\,
            I => \N__37445\
        );

    \I__7955\ : CascadeMux
    port map (
            O => \N__37449\,
            I => \N__37440\
        );

    \I__7954\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37437\
        );

    \I__7953\ : InMux
    port map (
            O => \N__37445\,
            I => \N__37432\
        );

    \I__7952\ : InMux
    port map (
            O => \N__37444\,
            I => \N__37432\
        );

    \I__7951\ : CascadeMux
    port map (
            O => \N__37443\,
            I => \N__37428\
        );

    \I__7950\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37424\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__37437\,
            I => \N__37421\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__37432\,
            I => \N__37418\
        );

    \I__7947\ : InMux
    port map (
            O => \N__37431\,
            I => \N__37413\
        );

    \I__7946\ : InMux
    port map (
            O => \N__37428\,
            I => \N__37413\
        );

    \I__7945\ : InMux
    port map (
            O => \N__37427\,
            I => \N__37410\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37405\
        );

    \I__7943\ : Span4Mux_v
    port map (
            O => \N__37421\,
            I => \N__37402\
        );

    \I__7942\ : Span4Mux_v
    port map (
            O => \N__37418\,
            I => \N__37399\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__37413\,
            I => \N__37394\
        );

    \I__7940\ : LocalMux
    port map (
            O => \N__37410\,
            I => \N__37394\
        );

    \I__7939\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37391\
        );

    \I__7938\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37388\
        );

    \I__7937\ : Span4Mux_v
    port map (
            O => \N__37405\,
            I => \N__37381\
        );

    \I__7936\ : Span4Mux_h
    port map (
            O => \N__37402\,
            I => \N__37381\
        );

    \I__7935\ : Span4Mux_h
    port map (
            O => \N__37399\,
            I => \N__37381\
        );

    \I__7934\ : Span4Mux_v
    port map (
            O => \N__37394\,
            I => \N__37376\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__37391\,
            I => \N__37376\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__37388\,
            I => \N__37373\
        );

    \I__7931\ : Span4Mux_v
    port map (
            O => \N__37381\,
            I => \N__37368\
        );

    \I__7930\ : Span4Mux_v
    port map (
            O => \N__37376\,
            I => \N__37368\
        );

    \I__7929\ : Odrv4
    port map (
            O => \N__37373\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__37368\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__7927\ : CascadeMux
    port map (
            O => \N__37363\,
            I => \N__37359\
        );

    \I__7926\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37356\
        );

    \I__7925\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37353\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__37356\,
            I => \N__37350\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__37353\,
            I => \N__37347\
        );

    \I__7922\ : Span4Mux_v
    port map (
            O => \N__37350\,
            I => \N__37344\
        );

    \I__7921\ : Span4Mux_v
    port map (
            O => \N__37347\,
            I => \N__37341\
        );

    \I__7920\ : Span4Mux_h
    port map (
            O => \N__37344\,
            I => \N__37338\
        );

    \I__7919\ : Sp12to4
    port map (
            O => \N__37341\,
            I => \N__37335\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__37338\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\
        );

    \I__7917\ : Odrv12
    port map (
            O => \N__37335\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\
        );

    \I__7916\ : InMux
    port map (
            O => \N__37330\,
            I => \N__37323\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37323\
        );

    \I__7914\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37318\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__37323\,
            I => \N__37314\
        );

    \I__7912\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37309\
        );

    \I__7911\ : InMux
    port map (
            O => \N__37321\,
            I => \N__37309\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__37318\,
            I => \N__37306\
        );

    \I__7909\ : InMux
    port map (
            O => \N__37317\,
            I => \N__37303\
        );

    \I__7908\ : Odrv12
    port map (
            O => \N__37314\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__37309\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__7906\ : Odrv4
    port map (
            O => \N__37306\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__37303\,
            I => \current_shift_inst.elapsed_time_ns_phase_1\
        );

    \I__7904\ : InMux
    port map (
            O => \N__37294\,
            I => \N__37290\
        );

    \I__7903\ : CascadeMux
    port map (
            O => \N__37293\,
            I => \N__37287\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__37290\,
            I => \N__37282\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37277\
        );

    \I__7900\ : InMux
    port map (
            O => \N__37286\,
            I => \N__37277\
        );

    \I__7899\ : InMux
    port map (
            O => \N__37285\,
            I => \N__37274\
        );

    \I__7898\ : Odrv12
    port map (
            O => \N__37282\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__37277\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__37274\,
            I => \current_shift_inst.elapsed_time_ns_phase_2\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37267\,
            I => \N__37264\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__37264\,
            I => \N__37261\
        );

    \I__7893\ : Odrv4
    port map (
            O => \N__37261\,
            I => \current_shift_inst.z_5_2\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37258\,
            I => \current_shift_inst.z_5_cry_1\
        );

    \I__7891\ : InMux
    port map (
            O => \N__37255\,
            I => \N__37252\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__37252\,
            I => \N__37249\
        );

    \I__7889\ : Odrv4
    port map (
            O => \N__37249\,
            I => \current_shift_inst.z_5_3\
        );

    \I__7888\ : InMux
    port map (
            O => \N__37246\,
            I => \current_shift_inst.z_5_cry_2\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__37243\,
            I => \N__37240\
        );

    \I__7886\ : InMux
    port map (
            O => \N__37240\,
            I => \N__37237\
        );

    \I__7885\ : LocalMux
    port map (
            O => \N__37237\,
            I => \N__37234\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__37234\,
            I => \current_shift_inst.z_5_4\
        );

    \I__7883\ : InMux
    port map (
            O => \N__37231\,
            I => \current_shift_inst.z_5_cry_3\
        );

    \I__7882\ : InMux
    port map (
            O => \N__37228\,
            I => \N__37225\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37225\,
            I => \N__37222\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__37222\,
            I => \current_shift_inst.z_5_5\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37219\,
            I => \current_shift_inst.z_5_cry_4\
        );

    \I__7878\ : CascadeMux
    port map (
            O => \N__37216\,
            I => \N__37213\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37213\,
            I => \N__37210\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__37210\,
            I => \N__37207\
        );

    \I__7875\ : Odrv4
    port map (
            O => \N__37207\,
            I => \current_shift_inst.z_5_6\
        );

    \I__7874\ : InMux
    port map (
            O => \N__37204\,
            I => \current_shift_inst.z_5_cry_5\
        );

    \I__7873\ : InMux
    port map (
            O => \N__37201\,
            I => \N__37198\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__37198\,
            I => \N__37195\
        );

    \I__7871\ : Odrv4
    port map (
            O => \N__37195\,
            I => \current_shift_inst.un4_control_input_axb_21\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37192\,
            I => \N__37189\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__37189\,
            I => \N__37186\
        );

    \I__7868\ : Span4Mux_h
    port map (
            O => \N__37186\,
            I => \N__37183\
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__37183\,
            I => \current_shift_inst.un4_control_input_axb_13\
        );

    \I__7866\ : InMux
    port map (
            O => \N__37180\,
            I => \N__37176\
        );

    \I__7865\ : InMux
    port map (
            O => \N__37179\,
            I => \N__37173\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__37176\,
            I => \N__37169\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__37173\,
            I => \N__37166\
        );

    \I__7862\ : InMux
    port map (
            O => \N__37172\,
            I => \N__37163\
        );

    \I__7861\ : Span4Mux_v
    port map (
            O => \N__37169\,
            I => \N__37158\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__37166\,
            I => \N__37158\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__37163\,
            I => measured_delay_tr_12
        );

    \I__7858\ : Odrv4
    port map (
            O => \N__37158\,
            I => measured_delay_tr_12
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__37153\,
            I => \N__37149\
        );

    \I__7856\ : InMux
    port map (
            O => \N__37152\,
            I => \N__37145\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37142\
        );

    \I__7854\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37139\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__37145\,
            I => \N__37134\
        );

    \I__7852\ : LocalMux
    port map (
            O => \N__37142\,
            I => \N__37134\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37139\,
            I => measured_delay_tr_13
        );

    \I__7850\ : Odrv12
    port map (
            O => \N__37134\,
            I => measured_delay_tr_13
        );

    \I__7849\ : InMux
    port map (
            O => \N__37129\,
            I => \N__37124\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37128\,
            I => \N__37121\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37118\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__37124\,
            I => \N__37113\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__37121\,
            I => \N__37113\
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__37118\,
            I => measured_delay_tr_11
        );

    \I__7843\ : Odrv12
    port map (
            O => \N__37113\,
            I => measured_delay_tr_11
        );

    \I__7842\ : InMux
    port map (
            O => \N__37108\,
            I => \N__37103\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37100\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37097\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__37103\,
            I => \N__37092\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__37100\,
            I => \N__37092\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__37097\,
            I => measured_delay_tr_10
        );

    \I__7836\ : Odrv12
    port map (
            O => \N__37092\,
            I => measured_delay_tr_10
        );

    \I__7835\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37084\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37084\,
            I => \current_shift_inst.un4_control_input_axb_30\
        );

    \I__7833\ : InMux
    port map (
            O => \N__37081\,
            I => \N__37078\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__37078\,
            I => \current_shift_inst.un4_control_input_axb_26\
        );

    \I__7831\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37072\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__37072\,
            I => \current_shift_inst.un4_control_input_axb_29\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37069\,
            I => \N__37066\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__37066\,
            I => \current_shift_inst.un4_control_input_axb_28\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37063\,
            I => \N__37060\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__37060\,
            I => \current_shift_inst.un4_control_input_axb_25\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__37057\,
            I => \N__37054\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37051\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__37051\,
            I => \N__37048\
        );

    \I__7822\ : Span4Mux_v
    port map (
            O => \N__37048\,
            I => \N__37045\
        );

    \I__7821\ : Odrv4
    port map (
            O => \N__37045\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__7820\ : CascadeMux
    port map (
            O => \N__37042\,
            I => \N__37039\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37039\,
            I => \N__37036\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__37036\,
            I => \N__37033\
        );

    \I__7817\ : Span4Mux_v
    port map (
            O => \N__37033\,
            I => \N__37030\
        );

    \I__7816\ : Odrv4
    port map (
            O => \N__37030\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__7815\ : CascadeMux
    port map (
            O => \N__37027\,
            I => \N__37024\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37024\,
            I => \N__37021\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37021\,
            I => \N__37018\
        );

    \I__7812\ : Span4Mux_v
    port map (
            O => \N__37018\,
            I => \N__37015\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__37015\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__37012\,
            I => \N__37006\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37011\,
            I => \N__37002\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37010\,
            I => \N__36993\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37009\,
            I => \N__36993\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37006\,
            I => \N__36993\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37005\,
            I => \N__36993\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__37002\,
            I => \N__36986\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36983\
        );

    \I__7802\ : InMux
    port map (
            O => \N__36992\,
            I => \N__36974\
        );

    \I__7801\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36974\
        );

    \I__7800\ : InMux
    port map (
            O => \N__36990\,
            I => \N__36974\
        );

    \I__7799\ : InMux
    port map (
            O => \N__36989\,
            I => \N__36974\
        );

    \I__7798\ : Span4Mux_v
    port map (
            O => \N__36986\,
            I => \N__36966\
        );

    \I__7797\ : Span4Mux_v
    port map (
            O => \N__36983\,
            I => \N__36966\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__36974\,
            I => \N__36966\
        );

    \I__7795\ : InMux
    port map (
            O => \N__36973\,
            I => \N__36963\
        );

    \I__7794\ : Span4Mux_v
    port map (
            O => \N__36966\,
            I => \N__36958\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__36963\,
            I => \N__36958\
        );

    \I__7792\ : Span4Mux_h
    port map (
            O => \N__36958\,
            I => \N__36955\
        );

    \I__7791\ : Odrv4
    port map (
            O => \N__36955\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__36952\,
            I => \N__36949\
        );

    \I__7789\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36946\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__36946\,
            I => \N__36943\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__36943\,
            I => \N__36940\
        );

    \I__7786\ : Span4Mux_v
    port map (
            O => \N__36940\,
            I => \N__36937\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__36937\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__7784\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36931\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__36931\,
            I => \current_shift_inst.un4_control_input_axb_12\
        );

    \I__7782\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36925\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__36925\,
            I => \current_shift_inst.un4_control_input_axb_19\
        );

    \I__7780\ : InMux
    port map (
            O => \N__36922\,
            I => \N__36919\
        );

    \I__7779\ : LocalMux
    port map (
            O => \N__36919\,
            I => \current_shift_inst.un4_control_input_axb_17\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__36916\,
            I => \N__36913\
        );

    \I__7777\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36910\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__36910\,
            I => \current_shift_inst.un4_control_input_axb_15\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__36907\,
            I => \N__36904\
        );

    \I__7774\ : InMux
    port map (
            O => \N__36904\,
            I => \N__36901\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__36901\,
            I => \current_shift_inst.un4_control_input_axb_16\
        );

    \I__7772\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36895\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__36895\,
            I => \current_shift_inst.un4_control_input_axb_18\
        );

    \I__7770\ : InMux
    port map (
            O => \N__36892\,
            I => \N__36889\
        );

    \I__7769\ : LocalMux
    port map (
            O => \N__36889\,
            I => \current_shift_inst.un4_control_input_axb_23\
        );

    \I__7768\ : InMux
    port map (
            O => \N__36886\,
            I => \N__36883\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__36883\,
            I => \current_shift_inst.un4_control_input_axb_27\
        );

    \I__7766\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36877\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__36877\,
            I => \current_shift_inst.un4_control_input_axb_20\
        );

    \I__7764\ : InMux
    port map (
            O => \N__36874\,
            I => \N__36871\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__36871\,
            I => \current_shift_inst.un4_control_input_axb_6\
        );

    \I__7762\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36865\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__36865\,
            I => \current_shift_inst.un4_control_input_axb_7\
        );

    \I__7760\ : InMux
    port map (
            O => \N__36862\,
            I => \N__36859\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__36859\,
            I => \current_shift_inst.un4_control_input_axb_8\
        );

    \I__7758\ : InMux
    port map (
            O => \N__36856\,
            I => \N__36853\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__36853\,
            I => \current_shift_inst.un4_control_input_axb_9\
        );

    \I__7756\ : InMux
    port map (
            O => \N__36850\,
            I => \N__36847\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__36847\,
            I => \current_shift_inst.un4_control_input_axb_10\
        );

    \I__7754\ : InMux
    port map (
            O => \N__36844\,
            I => \N__36841\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__36841\,
            I => \current_shift_inst.un4_control_input_axb_11\
        );

    \I__7752\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36835\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__36835\,
            I => \current_shift_inst.un4_control_input_axb_22\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__36832\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_\
        );

    \I__7749\ : InMux
    port map (
            O => \N__36829\,
            I => \N__36823\
        );

    \I__7748\ : InMux
    port map (
            O => \N__36828\,
            I => \N__36823\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__36823\,
            I => \N__36818\
        );

    \I__7746\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36815\
        );

    \I__7745\ : CascadeMux
    port map (
            O => \N__36821\,
            I => \N__36812\
        );

    \I__7744\ : Span4Mux_h
    port map (
            O => \N__36818\,
            I => \N__36808\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__36815\,
            I => \N__36805\
        );

    \I__7742\ : InMux
    port map (
            O => \N__36812\,
            I => \N__36802\
        );

    \I__7741\ : InMux
    port map (
            O => \N__36811\,
            I => \N__36799\
        );

    \I__7740\ : Span4Mux_v
    port map (
            O => \N__36808\,
            I => \N__36796\
        );

    \I__7739\ : Span4Mux_h
    port map (
            O => \N__36805\,
            I => \N__36793\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__36802\,
            I => measured_delay_tr_14
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__36799\,
            I => measured_delay_tr_14
        );

    \I__7736\ : Odrv4
    port map (
            O => \N__36796\,
            I => measured_delay_tr_14
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__36793\,
            I => measured_delay_tr_14
        );

    \I__7734\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36781\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__36781\,
            I => \current_shift_inst.un4_control_input_axb_4\
        );

    \I__7732\ : InMux
    port map (
            O => \N__36778\,
            I => \N__36775\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__36775\,
            I => \current_shift_inst.un4_control_input_axb_5\
        );

    \I__7730\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36769\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__36769\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__36766\,
            I => \N__36763\
        );

    \I__7727\ : InMux
    port map (
            O => \N__36763\,
            I => \N__36760\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__36760\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__7725\ : InMux
    port map (
            O => \N__36757\,
            I => \N__36754\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36754\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__7723\ : CascadeMux
    port map (
            O => \N__36751\,
            I => \N__36748\
        );

    \I__7722\ : InMux
    port map (
            O => \N__36748\,
            I => \N__36745\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36745\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__7720\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36739\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__36739\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__7718\ : InMux
    port map (
            O => \N__36736\,
            I => \N__36733\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__36733\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__7716\ : CascadeMux
    port map (
            O => \N__36730\,
            I => \N__36727\
        );

    \I__7715\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36724\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__36724\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__7713\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36718\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__36718\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__7711\ : CascadeMux
    port map (
            O => \N__36715\,
            I => \N__36712\
        );

    \I__7710\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36709\
        );

    \I__7709\ : LocalMux
    port map (
            O => \N__36709\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36706\,
            I => \N__36703\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__36703\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__7706\ : CascadeMux
    port map (
            O => \N__36700\,
            I => \N__36697\
        );

    \I__7705\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36694\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__36694\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__36691\,
            I => \N__36688\
        );

    \I__7702\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36685\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__36685\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__7700\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36679\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__36679\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__36676\,
            I => \N__36673\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36673\,
            I => \N__36670\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__36670\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__7695\ : InMux
    port map (
            O => \N__36667\,
            I => \N__36643\
        );

    \I__7694\ : InMux
    port map (
            O => \N__36666\,
            I => \N__36630\
        );

    \I__7693\ : InMux
    port map (
            O => \N__36665\,
            I => \N__36630\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36630\
        );

    \I__7691\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36630\
        );

    \I__7690\ : InMux
    port map (
            O => \N__36662\,
            I => \N__36630\
        );

    \I__7689\ : InMux
    port map (
            O => \N__36661\,
            I => \N__36630\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36660\,
            I => \N__36615\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36659\,
            I => \N__36615\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36658\,
            I => \N__36615\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36615\
        );

    \I__7684\ : InMux
    port map (
            O => \N__36656\,
            I => \N__36615\
        );

    \I__7683\ : InMux
    port map (
            O => \N__36655\,
            I => \N__36615\
        );

    \I__7682\ : InMux
    port map (
            O => \N__36654\,
            I => \N__36615\
        );

    \I__7681\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36596\
        );

    \I__7680\ : InMux
    port map (
            O => \N__36652\,
            I => \N__36596\
        );

    \I__7679\ : InMux
    port map (
            O => \N__36651\,
            I => \N__36596\
        );

    \I__7678\ : InMux
    port map (
            O => \N__36650\,
            I => \N__36596\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36596\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36648\,
            I => \N__36596\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36647\,
            I => \N__36596\
        );

    \I__7674\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36593\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36588\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__36630\,
            I => \N__36588\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__36615\,
            I => \N__36581\
        );

    \I__7670\ : InMux
    port map (
            O => \N__36614\,
            I => \N__36572\
        );

    \I__7669\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36572\
        );

    \I__7668\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36572\
        );

    \I__7667\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36572\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__36596\,
            I => \N__36567\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__36593\,
            I => \N__36567\
        );

    \I__7664\ : Span4Mux_v
    port map (
            O => \N__36588\,
            I => \N__36558\
        );

    \I__7663\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36549\
        );

    \I__7662\ : InMux
    port map (
            O => \N__36586\,
            I => \N__36549\
        );

    \I__7661\ : InMux
    port map (
            O => \N__36585\,
            I => \N__36549\
        );

    \I__7660\ : InMux
    port map (
            O => \N__36584\,
            I => \N__36549\
        );

    \I__7659\ : Span4Mux_v
    port map (
            O => \N__36581\,
            I => \N__36544\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__36572\,
            I => \N__36544\
        );

    \I__7657\ : Span4Mux_h
    port map (
            O => \N__36567\,
            I => \N__36541\
        );

    \I__7656\ : InMux
    port map (
            O => \N__36566\,
            I => \N__36534\
        );

    \I__7655\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36534\
        );

    \I__7654\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36534\
        );

    \I__7653\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36527\
        );

    \I__7652\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36527\
        );

    \I__7651\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36527\
        );

    \I__7650\ : Sp12to4
    port map (
            O => \N__36558\,
            I => \N__36520\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36520\
        );

    \I__7648\ : Span4Mux_h
    port map (
            O => \N__36544\,
            I => \N__36517\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__36541\,
            I => \N__36510\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__36534\,
            I => \N__36510\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__36527\,
            I => \N__36510\
        );

    \I__7644\ : InMux
    port map (
            O => \N__36526\,
            I => \N__36505\
        );

    \I__7643\ : InMux
    port map (
            O => \N__36525\,
            I => \N__36505\
        );

    \I__7642\ : Odrv12
    port map (
            O => \N__36520\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7641\ : Odrv4
    port map (
            O => \N__36517\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7640\ : Odrv4
    port map (
            O => \N__36510\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__36505\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt31_0\
        );

    \I__7638\ : InMux
    port map (
            O => \N__36496\,
            I => \N__36492\
        );

    \I__7637\ : CascadeMux
    port map (
            O => \N__36495\,
            I => \N__36487\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__36492\,
            I => \N__36484\
        );

    \I__7635\ : InMux
    port map (
            O => \N__36491\,
            I => \N__36481\
        );

    \I__7634\ : InMux
    port map (
            O => \N__36490\,
            I => \N__36478\
        );

    \I__7633\ : InMux
    port map (
            O => \N__36487\,
            I => \N__36474\
        );

    \I__7632\ : Span4Mux_h
    port map (
            O => \N__36484\,
            I => \N__36471\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__36481\,
            I => \N__36468\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__36478\,
            I => \N__36465\
        );

    \I__7629\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36462\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__36474\,
            I => measured_delay_hc_8
        );

    \I__7627\ : Odrv4
    port map (
            O => \N__36471\,
            I => measured_delay_hc_8
        );

    \I__7626\ : Odrv12
    port map (
            O => \N__36468\,
            I => measured_delay_hc_8
        );

    \I__7625\ : Odrv4
    port map (
            O => \N__36465\,
            I => measured_delay_hc_8
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__36462\,
            I => measured_delay_hc_8
        );

    \I__7623\ : CascadeMux
    port map (
            O => \N__36451\,
            I => \N__36446\
        );

    \I__7622\ : CascadeMux
    port map (
            O => \N__36450\,
            I => \N__36434\
        );

    \I__7621\ : CascadeMux
    port map (
            O => \N__36449\,
            I => \N__36431\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36446\,
            I => \N__36422\
        );

    \I__7619\ : InMux
    port map (
            O => \N__36445\,
            I => \N__36422\
        );

    \I__7618\ : InMux
    port map (
            O => \N__36444\,
            I => \N__36422\
        );

    \I__7617\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36422\
        );

    \I__7616\ : CascadeMux
    port map (
            O => \N__36442\,
            I => \N__36414\
        );

    \I__7615\ : InMux
    port map (
            O => \N__36441\,
            I => \N__36399\
        );

    \I__7614\ : InMux
    port map (
            O => \N__36440\,
            I => \N__36399\
        );

    \I__7613\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36399\
        );

    \I__7612\ : InMux
    port map (
            O => \N__36438\,
            I => \N__36399\
        );

    \I__7611\ : InMux
    port map (
            O => \N__36437\,
            I => \N__36399\
        );

    \I__7610\ : InMux
    port map (
            O => \N__36434\,
            I => \N__36399\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36399\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__36422\,
            I => \N__36393\
        );

    \I__7607\ : InMux
    port map (
            O => \N__36421\,
            I => \N__36386\
        );

    \I__7606\ : InMux
    port map (
            O => \N__36420\,
            I => \N__36386\
        );

    \I__7605\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36386\
        );

    \I__7604\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36379\
        );

    \I__7603\ : InMux
    port map (
            O => \N__36417\,
            I => \N__36379\
        );

    \I__7602\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36379\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__36399\,
            I => \N__36376\
        );

    \I__7600\ : InMux
    port map (
            O => \N__36398\,
            I => \N__36369\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36369\
        );

    \I__7598\ : InMux
    port map (
            O => \N__36396\,
            I => \N__36369\
        );

    \I__7597\ : Span4Mux_h
    port map (
            O => \N__36393\,
            I => \N__36362\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__36386\,
            I => \N__36362\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__36379\,
            I => \N__36354\
        );

    \I__7594\ : Span4Mux_h
    port map (
            O => \N__36376\,
            I => \N__36349\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__36369\,
            I => \N__36349\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__36368\,
            I => \N__36345\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__36367\,
            I => \N__36341\
        );

    \I__7590\ : Span4Mux_v
    port map (
            O => \N__36362\,
            I => \N__36336\
        );

    \I__7589\ : CascadeMux
    port map (
            O => \N__36361\,
            I => \N__36332\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__36360\,
            I => \N__36329\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__36359\,
            I => \N__36326\
        );

    \I__7586\ : CascadeMux
    port map (
            O => \N__36358\,
            I => \N__36322\
        );

    \I__7585\ : CascadeMux
    port map (
            O => \N__36357\,
            I => \N__36311\
        );

    \I__7584\ : Span4Mux_v
    port map (
            O => \N__36354\,
            I => \N__36306\
        );

    \I__7583\ : Span4Mux_h
    port map (
            O => \N__36349\,
            I => \N__36306\
        );

    \I__7582\ : InMux
    port map (
            O => \N__36348\,
            I => \N__36295\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36295\
        );

    \I__7580\ : InMux
    port map (
            O => \N__36344\,
            I => \N__36295\
        );

    \I__7579\ : InMux
    port map (
            O => \N__36341\,
            I => \N__36295\
        );

    \I__7578\ : InMux
    port map (
            O => \N__36340\,
            I => \N__36295\
        );

    \I__7577\ : InMux
    port map (
            O => \N__36339\,
            I => \N__36292\
        );

    \I__7576\ : Span4Mux_h
    port map (
            O => \N__36336\,
            I => \N__36289\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36335\,
            I => \N__36286\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36271\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36329\,
            I => \N__36271\
        );

    \I__7572\ : InMux
    port map (
            O => \N__36326\,
            I => \N__36271\
        );

    \I__7571\ : InMux
    port map (
            O => \N__36325\,
            I => \N__36271\
        );

    \I__7570\ : InMux
    port map (
            O => \N__36322\,
            I => \N__36271\
        );

    \I__7569\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36271\
        );

    \I__7568\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36271\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36268\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36255\
        );

    \I__7565\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36255\
        );

    \I__7564\ : InMux
    port map (
            O => \N__36316\,
            I => \N__36255\
        );

    \I__7563\ : InMux
    port map (
            O => \N__36315\,
            I => \N__36255\
        );

    \I__7562\ : InMux
    port map (
            O => \N__36314\,
            I => \N__36255\
        );

    \I__7561\ : InMux
    port map (
            O => \N__36311\,
            I => \N__36255\
        );

    \I__7560\ : Span4Mux_h
    port map (
            O => \N__36306\,
            I => \N__36250\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__36295\,
            I => \N__36250\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36292\,
            I => measured_delay_hc_31
        );

    \I__7557\ : Odrv4
    port map (
            O => \N__36289\,
            I => measured_delay_hc_31
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__36286\,
            I => measured_delay_hc_31
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__36271\,
            I => measured_delay_hc_31
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__36268\,
            I => measured_delay_hc_31
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__36255\,
            I => measured_delay_hc_31
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__36250\,
            I => measured_delay_hc_31
        );

    \I__7551\ : CascadeMux
    port map (
            O => \N__36235\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__7550\ : CEMux
    port map (
            O => \N__36232\,
            I => \N__36228\
        );

    \I__7549\ : CEMux
    port map (
            O => \N__36231\,
            I => \N__36223\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__36228\,
            I => \N__36219\
        );

    \I__7547\ : CEMux
    port map (
            O => \N__36227\,
            I => \N__36216\
        );

    \I__7546\ : CEMux
    port map (
            O => \N__36226\,
            I => \N__36213\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36223\,
            I => \N__36210\
        );

    \I__7544\ : CEMux
    port map (
            O => \N__36222\,
            I => \N__36207\
        );

    \I__7543\ : Span4Mux_v
    port map (
            O => \N__36219\,
            I => \N__36202\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__36216\,
            I => \N__36202\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__36213\,
            I => \N__36199\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__36210\,
            I => \N__36196\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__36207\,
            I => \N__36193\
        );

    \I__7538\ : Span4Mux_h
    port map (
            O => \N__36202\,
            I => \N__36190\
        );

    \I__7537\ : Span4Mux_v
    port map (
            O => \N__36199\,
            I => \N__36185\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__36196\,
            I => \N__36185\
        );

    \I__7535\ : Odrv12
    port map (
            O => \N__36193\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__36190\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__36185\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36178\,
            I => \N__36175\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__36175\,
            I => \N__36172\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__36172\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36169\,
            I => \N__36166\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__36166\,
            I => \N__36163\
        );

    \I__7527\ : Odrv4
    port map (
            O => \N__36163\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__7526\ : CascadeMux
    port map (
            O => \N__36160\,
            I => \N__36157\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36157\,
            I => \N__36154\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36154\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36146\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36150\,
            I => \N__36143\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36149\,
            I => \N__36140\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__36146\,
            I => \N__36136\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__36143\,
            I => \N__36133\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36130\
        );

    \I__7517\ : CascadeMux
    port map (
            O => \N__36139\,
            I => \N__36126\
        );

    \I__7516\ : Span4Mux_h
    port map (
            O => \N__36136\,
            I => \N__36123\
        );

    \I__7515\ : Span4Mux_v
    port map (
            O => \N__36133\,
            I => \N__36120\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36130\,
            I => \N__36117\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36114\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36111\
        );

    \I__7511\ : Span4Mux_h
    port map (
            O => \N__36123\,
            I => \N__36108\
        );

    \I__7510\ : Span4Mux_h
    port map (
            O => \N__36120\,
            I => \N__36101\
        );

    \I__7509\ : Span4Mux_v
    port map (
            O => \N__36117\,
            I => \N__36101\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__36114\,
            I => \N__36101\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__36111\,
            I => measured_delay_hc_5
        );

    \I__7506\ : Odrv4
    port map (
            O => \N__36108\,
            I => measured_delay_hc_5
        );

    \I__7505\ : Odrv4
    port map (
            O => \N__36101\,
            I => measured_delay_hc_5
        );

    \I__7504\ : CascadeMux
    port map (
            O => \N__36094\,
            I => \N__36091\
        );

    \I__7503\ : InMux
    port map (
            O => \N__36091\,
            I => \N__36088\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__36088\,
            I => \N__36082\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36087\,
            I => \N__36079\
        );

    \I__7500\ : CascadeMux
    port map (
            O => \N__36086\,
            I => \N__36076\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36073\
        );

    \I__7498\ : Span4Mux_h
    port map (
            O => \N__36082\,
            I => \N__36070\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36079\,
            I => \N__36067\
        );

    \I__7496\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36064\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__36073\,
            I => \N__36060\
        );

    \I__7494\ : Span4Mux_h
    port map (
            O => \N__36070\,
            I => \N__36055\
        );

    \I__7493\ : Span4Mux_h
    port map (
            O => \N__36067\,
            I => \N__36055\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__36064\,
            I => \N__36052\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36063\,
            I => \N__36049\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__36060\,
            I => \N__36046\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__36055\,
            I => \N__36043\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__36052\,
            I => \N__36040\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36049\,
            I => measured_delay_hc_3
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__36046\,
            I => measured_delay_hc_3
        );

    \I__7485\ : Odrv4
    port map (
            O => \N__36043\,
            I => measured_delay_hc_3
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__36040\,
            I => measured_delay_hc_3
        );

    \I__7483\ : InMux
    port map (
            O => \N__36031\,
            I => \N__36028\
        );

    \I__7482\ : LocalMux
    port map (
            O => \N__36028\,
            I => \N__36024\
        );

    \I__7481\ : InMux
    port map (
            O => \N__36027\,
            I => \N__36021\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__36024\,
            I => \N__36015\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__36012\
        );

    \I__7478\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36009\
        );

    \I__7477\ : CascadeMux
    port map (
            O => \N__36019\,
            I => \N__36006\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36018\,
            I => \N__36003\
        );

    \I__7475\ : Span4Mux_h
    port map (
            O => \N__36015\,
            I => \N__35996\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__36012\,
            I => \N__35996\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__36009\,
            I => \N__35996\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35993\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__36003\,
            I => measured_delay_hc_13
        );

    \I__7470\ : Odrv4
    port map (
            O => \N__35996\,
            I => measured_delay_hc_13
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__35993\,
            I => measured_delay_hc_13
        );

    \I__7468\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35980\
        );

    \I__7467\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35977\
        );

    \I__7466\ : CascadeMux
    port map (
            O => \N__35984\,
            I => \N__35974\
        );

    \I__7465\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35971\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__35980\,
            I => \N__35968\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__35977\,
            I => \N__35963\
        );

    \I__7462\ : InMux
    port map (
            O => \N__35974\,
            I => \N__35960\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__35971\,
            I => \N__35957\
        );

    \I__7460\ : Span4Mux_v
    port map (
            O => \N__35968\,
            I => \N__35954\
        );

    \I__7459\ : InMux
    port map (
            O => \N__35967\,
            I => \N__35951\
        );

    \I__7458\ : InMux
    port map (
            O => \N__35966\,
            I => \N__35948\
        );

    \I__7457\ : Span4Mux_h
    port map (
            O => \N__35963\,
            I => \N__35945\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__35960\,
            I => measured_delay_hc_9
        );

    \I__7455\ : Odrv12
    port map (
            O => \N__35957\,
            I => measured_delay_hc_9
        );

    \I__7454\ : Odrv4
    port map (
            O => \N__35954\,
            I => measured_delay_hc_9
        );

    \I__7453\ : LocalMux
    port map (
            O => \N__35951\,
            I => measured_delay_hc_9
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__35948\,
            I => measured_delay_hc_9
        );

    \I__7451\ : Odrv4
    port map (
            O => \N__35945\,
            I => measured_delay_hc_9
        );

    \I__7450\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35927\
        );

    \I__7449\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35924\
        );

    \I__7448\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35920\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__35927\,
            I => \N__35917\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__35924\,
            I => \N__35914\
        );

    \I__7445\ : InMux
    port map (
            O => \N__35923\,
            I => \N__35911\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__35920\,
            I => \N__35905\
        );

    \I__7443\ : Span4Mux_h
    port map (
            O => \N__35917\,
            I => \N__35905\
        );

    \I__7442\ : Span4Mux_h
    port map (
            O => \N__35914\,
            I => \N__35900\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__35911\,
            I => \N__35900\
        );

    \I__7440\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35897\
        );

    \I__7439\ : Odrv4
    port map (
            O => \N__35905\,
            I => measured_delay_hc_10
        );

    \I__7438\ : Odrv4
    port map (
            O => \N__35900\,
            I => measured_delay_hc_10
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__35897\,
            I => measured_delay_hc_10
        );

    \I__7436\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35885\
        );

    \I__7435\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35882\
        );

    \I__7434\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35878\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__35885\,
            I => \N__35875\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__35882\,
            I => \N__35872\
        );

    \I__7431\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35869\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35863\
        );

    \I__7429\ : Span4Mux_h
    port map (
            O => \N__35875\,
            I => \N__35863\
        );

    \I__7428\ : Span4Mux_h
    port map (
            O => \N__35872\,
            I => \N__35858\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__35869\,
            I => \N__35858\
        );

    \I__7426\ : InMux
    port map (
            O => \N__35868\,
            I => \N__35855\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__35863\,
            I => measured_delay_hc_11
        );

    \I__7424\ : Odrv4
    port map (
            O => \N__35858\,
            I => measured_delay_hc_11
        );

    \I__7423\ : LocalMux
    port map (
            O => \N__35855\,
            I => measured_delay_hc_11
        );

    \I__7422\ : CascadeMux
    port map (
            O => \N__35848\,
            I => \N__35845\
        );

    \I__7421\ : InMux
    port map (
            O => \N__35845\,
            I => \N__35842\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__35842\,
            I => \N__35838\
        );

    \I__7419\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35834\
        );

    \I__7418\ : Span4Mux_v
    port map (
            O => \N__35838\,
            I => \N__35831\
        );

    \I__7417\ : InMux
    port map (
            O => \N__35837\,
            I => \N__35828\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35824\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__35831\,
            I => \N__35819\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__35828\,
            I => \N__35819\
        );

    \I__7413\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35816\
        );

    \I__7412\ : Span4Mux_h
    port map (
            O => \N__35824\,
            I => \N__35813\
        );

    \I__7411\ : Span4Mux_h
    port map (
            O => \N__35819\,
            I => \N__35810\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__35816\,
            I => measured_delay_hc_0
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__35813\,
            I => measured_delay_hc_0
        );

    \I__7408\ : Odrv4
    port map (
            O => \N__35810\,
            I => measured_delay_hc_0
        );

    \I__7407\ : CascadeMux
    port map (
            O => \N__35803\,
            I => \N__35798\
        );

    \I__7406\ : CascadeMux
    port map (
            O => \N__35802\,
            I => \N__35795\
        );

    \I__7405\ : CascadeMux
    port map (
            O => \N__35801\,
            I => \N__35792\
        );

    \I__7404\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35781\
        );

    \I__7403\ : InMux
    port map (
            O => \N__35795\,
            I => \N__35781\
        );

    \I__7402\ : InMux
    port map (
            O => \N__35792\,
            I => \N__35781\
        );

    \I__7401\ : InMux
    port map (
            O => \N__35791\,
            I => \N__35781\
        );

    \I__7400\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35770\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__35781\,
            I => \N__35766\
        );

    \I__7398\ : InMux
    port map (
            O => \N__35780\,
            I => \N__35759\
        );

    \I__7397\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35759\
        );

    \I__7396\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35759\
        );

    \I__7395\ : InMux
    port map (
            O => \N__35777\,
            I => \N__35748\
        );

    \I__7394\ : InMux
    port map (
            O => \N__35776\,
            I => \N__35748\
        );

    \I__7393\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35748\
        );

    \I__7392\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35748\
        );

    \I__7391\ : InMux
    port map (
            O => \N__35773\,
            I => \N__35748\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__35770\,
            I => \N__35745\
        );

    \I__7389\ : InMux
    port map (
            O => \N__35769\,
            I => \N__35742\
        );

    \I__7388\ : Span4Mux_v
    port map (
            O => \N__35766\,
            I => \N__35737\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35759\,
            I => \N__35737\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__35748\,
            I => \N__35734\
        );

    \I__7385\ : Span4Mux_v
    port map (
            O => \N__35745\,
            I => \N__35729\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35742\,
            I => \N__35729\
        );

    \I__7383\ : Span4Mux_h
    port map (
            O => \N__35737\,
            I => \N__35726\
        );

    \I__7382\ : Span4Mux_h
    port map (
            O => \N__35734\,
            I => \N__35723\
        );

    \I__7381\ : Span4Mux_h
    port map (
            O => \N__35729\,
            I => \N__35720\
        );

    \I__7380\ : Odrv4
    port map (
            O => \N__35726\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__7379\ : Odrv4
    port map (
            O => \N__35723\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__7378\ : Odrv4
    port map (
            O => \N__35720\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35713\,
            I => \N__35710\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__35710\,
            I => \N__35705\
        );

    \I__7375\ : CascadeMux
    port map (
            O => \N__35709\,
            I => \N__35701\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35698\
        );

    \I__7373\ : Span4Mux_h
    port map (
            O => \N__35705\,
            I => \N__35695\
        );

    \I__7372\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35692\
        );

    \I__7371\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35688\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35685\
        );

    \I__7369\ : Span4Mux_h
    port map (
            O => \N__35695\,
            I => \N__35680\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__35692\,
            I => \N__35680\
        );

    \I__7367\ : InMux
    port map (
            O => \N__35691\,
            I => \N__35677\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__35688\,
            I => measured_delay_hc_1
        );

    \I__7365\ : Odrv12
    port map (
            O => \N__35685\,
            I => measured_delay_hc_1
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__35680\,
            I => measured_delay_hc_1
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__35677\,
            I => measured_delay_hc_1
        );

    \I__7362\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35665\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35659\
        );

    \I__7360\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35655\
        );

    \I__7359\ : CascadeMux
    port map (
            O => \N__35663\,
            I => \N__35652\
        );

    \I__7358\ : InMux
    port map (
            O => \N__35662\,
            I => \N__35649\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__35659\,
            I => \N__35646\
        );

    \I__7356\ : InMux
    port map (
            O => \N__35658\,
            I => \N__35643\
        );

    \I__7355\ : LocalMux
    port map (
            O => \N__35655\,
            I => \N__35640\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35637\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__35649\,
            I => \N__35634\
        );

    \I__7352\ : Span4Mux_h
    port map (
            O => \N__35646\,
            I => \N__35631\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__35643\,
            I => \N__35628\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__35640\,
            I => \N__35625\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__35637\,
            I => measured_delay_hc_15
        );

    \I__7348\ : Odrv12
    port map (
            O => \N__35634\,
            I => measured_delay_hc_15
        );

    \I__7347\ : Odrv4
    port map (
            O => \N__35631\,
            I => measured_delay_hc_15
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__35628\,
            I => measured_delay_hc_15
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__35625\,
            I => measured_delay_hc_15
        );

    \I__7344\ : InMux
    port map (
            O => \N__35614\,
            I => \current_shift_inst.timer_phase.counter_cry_26\
        );

    \I__7343\ : InMux
    port map (
            O => \N__35611\,
            I => \current_shift_inst.timer_phase.counter_cry_27\
        );

    \I__7342\ : InMux
    port map (
            O => \N__35608\,
            I => \N__35570\
        );

    \I__7341\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35570\
        );

    \I__7340\ : InMux
    port map (
            O => \N__35606\,
            I => \N__35570\
        );

    \I__7339\ : InMux
    port map (
            O => \N__35605\,
            I => \N__35570\
        );

    \I__7338\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35561\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35561\
        );

    \I__7336\ : InMux
    port map (
            O => \N__35602\,
            I => \N__35561\
        );

    \I__7335\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35561\
        );

    \I__7334\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35556\
        );

    \I__7333\ : InMux
    port map (
            O => \N__35599\,
            I => \N__35556\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35598\,
            I => \N__35547\
        );

    \I__7331\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35547\
        );

    \I__7330\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35547\
        );

    \I__7329\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35547\
        );

    \I__7328\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35538\
        );

    \I__7327\ : InMux
    port map (
            O => \N__35593\,
            I => \N__35538\
        );

    \I__7326\ : InMux
    port map (
            O => \N__35592\,
            I => \N__35538\
        );

    \I__7325\ : InMux
    port map (
            O => \N__35591\,
            I => \N__35538\
        );

    \I__7324\ : InMux
    port map (
            O => \N__35590\,
            I => \N__35529\
        );

    \I__7323\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35529\
        );

    \I__7322\ : InMux
    port map (
            O => \N__35588\,
            I => \N__35529\
        );

    \I__7321\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35529\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35520\
        );

    \I__7319\ : InMux
    port map (
            O => \N__35585\,
            I => \N__35520\
        );

    \I__7318\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35520\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35520\
        );

    \I__7316\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35511\
        );

    \I__7315\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35511\
        );

    \I__7314\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35511\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35579\,
            I => \N__35511\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35506\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__35561\,
            I => \N__35506\
        );

    \I__7310\ : LocalMux
    port map (
            O => \N__35556\,
            I => \N__35497\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__35547\,
            I => \N__35497\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__35538\,
            I => \N__35497\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__35529\,
            I => \N__35497\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35488\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__35511\,
            I => \N__35488\
        );

    \I__7304\ : Span4Mux_v
    port map (
            O => \N__35506\,
            I => \N__35488\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__35497\,
            I => \N__35488\
        );

    \I__7302\ : Odrv4
    port map (
            O => \N__35488\,
            I => \current_shift_inst.timer_phase.running_i\
        );

    \I__7301\ : InMux
    port map (
            O => \N__35485\,
            I => \current_shift_inst.timer_phase.counter_cry_28\
        );

    \I__7300\ : CEMux
    port map (
            O => \N__35482\,
            I => \N__35477\
        );

    \I__7299\ : CEMux
    port map (
            O => \N__35481\,
            I => \N__35473\
        );

    \I__7298\ : CEMux
    port map (
            O => \N__35480\,
            I => \N__35470\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__35477\,
            I => \N__35467\
        );

    \I__7296\ : CEMux
    port map (
            O => \N__35476\,
            I => \N__35464\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__35473\,
            I => \N__35459\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35459\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__35467\,
            I => \N__35454\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__35464\,
            I => \N__35454\
        );

    \I__7291\ : Span4Mux_v
    port map (
            O => \N__35459\,
            I => \N__35451\
        );

    \I__7290\ : Span4Mux_v
    port map (
            O => \N__35454\,
            I => \N__35446\
        );

    \I__7289\ : Span4Mux_h
    port map (
            O => \N__35451\,
            I => \N__35446\
        );

    \I__7288\ : Odrv4
    port map (
            O => \N__35446\,
            I => \current_shift_inst.timer_phase.N_192_i\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35440\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__35440\,
            I => \N__35437\
        );

    \I__7285\ : Odrv12
    port map (
            O => \N__35437\,
            I => delay_tr_input_c
        );

    \I__7284\ : InMux
    port map (
            O => \N__35434\,
            I => \N__35431\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__35431\,
            I => delay_tr_d1
        );

    \I__7282\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35425\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__35425\,
            I => \N__35420\
        );

    \I__7280\ : InMux
    port map (
            O => \N__35424\,
            I => \N__35417\
        );

    \I__7279\ : CascadeMux
    port map (
            O => \N__35423\,
            I => \N__35413\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__35420\,
            I => \N__35410\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__35417\,
            I => \N__35407\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35404\
        );

    \I__7275\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35400\
        );

    \I__7274\ : Span4Mux_h
    port map (
            O => \N__35410\,
            I => \N__35397\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__35407\,
            I => \N__35392\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__35404\,
            I => \N__35392\
        );

    \I__7271\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35389\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__35400\,
            I => measured_delay_hc_7
        );

    \I__7269\ : Odrv4
    port map (
            O => \N__35397\,
            I => measured_delay_hc_7
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__35392\,
            I => measured_delay_hc_7
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__35389\,
            I => measured_delay_hc_7
        );

    \I__7266\ : CascadeMux
    port map (
            O => \N__35380\,
            I => \N__35375\
        );

    \I__7265\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35371\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__35378\,
            I => \N__35367\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35364\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35374\,
            I => \N__35361\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__35371\,
            I => \N__35358\
        );

    \I__7260\ : InMux
    port map (
            O => \N__35370\,
            I => \N__35355\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35367\,
            I => \N__35352\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__35364\,
            I => \N__35349\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__35361\,
            I => \N__35346\
        );

    \I__7256\ : Span4Mux_v
    port map (
            O => \N__35358\,
            I => \N__35341\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__35355\,
            I => \N__35341\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__35352\,
            I => \N__35336\
        );

    \I__7253\ : Span4Mux_v
    port map (
            O => \N__35349\,
            I => \N__35336\
        );

    \I__7252\ : Span12Mux_h
    port map (
            O => \N__35346\,
            I => \N__35333\
        );

    \I__7251\ : Span4Mux_h
    port map (
            O => \N__35341\,
            I => \N__35330\
        );

    \I__7250\ : Odrv4
    port map (
            O => \N__35336\,
            I => measured_delay_hc_2
        );

    \I__7249\ : Odrv12
    port map (
            O => \N__35333\,
            I => measured_delay_hc_2
        );

    \I__7248\ : Odrv4
    port map (
            O => \N__35330\,
            I => measured_delay_hc_2
        );

    \I__7247\ : InMux
    port map (
            O => \N__35323\,
            I => \N__35320\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__35320\,
            I => \N__35316\
        );

    \I__7245\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35310\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__35316\,
            I => \N__35307\
        );

    \I__7243\ : InMux
    port map (
            O => \N__35315\,
            I => \N__35304\
        );

    \I__7242\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35301\
        );

    \I__7241\ : CascadeMux
    port map (
            O => \N__35313\,
            I => \N__35298\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__35310\,
            I => \N__35295\
        );

    \I__7239\ : Sp12to4
    port map (
            O => \N__35307\,
            I => \N__35290\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__35304\,
            I => \N__35290\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__35301\,
            I => \N__35287\
        );

    \I__7236\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35284\
        );

    \I__7235\ : Span12Mux_h
    port map (
            O => \N__35295\,
            I => \N__35281\
        );

    \I__7234\ : Span12Mux_h
    port map (
            O => \N__35290\,
            I => \N__35278\
        );

    \I__7233\ : Span4Mux_h
    port map (
            O => \N__35287\,
            I => \N__35275\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__35284\,
            I => measured_delay_hc_6
        );

    \I__7231\ : Odrv12
    port map (
            O => \N__35281\,
            I => measured_delay_hc_6
        );

    \I__7230\ : Odrv12
    port map (
            O => \N__35278\,
            I => measured_delay_hc_6
        );

    \I__7229\ : Odrv4
    port map (
            O => \N__35275\,
            I => measured_delay_hc_6
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__35266\,
            I => \N__35262\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35265\,
            I => \N__35259\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35262\,
            I => \N__35256\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__35259\,
            I => \N__35251\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__35256\,
            I => \N__35248\
        );

    \I__7223\ : InMux
    port map (
            O => \N__35255\,
            I => \N__35245\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35254\,
            I => \N__35241\
        );

    \I__7221\ : Span4Mux_v
    port map (
            O => \N__35251\,
            I => \N__35238\
        );

    \I__7220\ : Span4Mux_h
    port map (
            O => \N__35248\,
            I => \N__35235\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__35245\,
            I => \N__35232\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35244\,
            I => \N__35229\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__35241\,
            I => \N__35226\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__35238\,
            I => \N__35219\
        );

    \I__7215\ : Span4Mux_v
    port map (
            O => \N__35235\,
            I => \N__35219\
        );

    \I__7214\ : Span4Mux_v
    port map (
            O => \N__35232\,
            I => \N__35219\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35229\,
            I => measured_delay_hc_4
        );

    \I__7212\ : Odrv4
    port map (
            O => \N__35226\,
            I => measured_delay_hc_4
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__35219\,
            I => measured_delay_hc_4
        );

    \I__7210\ : InMux
    port map (
            O => \N__35212\,
            I => \current_shift_inst.timer_phase.counter_cry_17\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35209\,
            I => \current_shift_inst.timer_phase.counter_cry_18\
        );

    \I__7208\ : InMux
    port map (
            O => \N__35206\,
            I => \current_shift_inst.timer_phase.counter_cry_19\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35203\,
            I => \current_shift_inst.timer_phase.counter_cry_20\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35200\,
            I => \current_shift_inst.timer_phase.counter_cry_21\
        );

    \I__7205\ : InMux
    port map (
            O => \N__35197\,
            I => \current_shift_inst.timer_phase.counter_cry_22\
        );

    \I__7204\ : InMux
    port map (
            O => \N__35194\,
            I => \bfn_14_25_0_\
        );

    \I__7203\ : InMux
    port map (
            O => \N__35191\,
            I => \current_shift_inst.timer_phase.counter_cry_24\
        );

    \I__7202\ : InMux
    port map (
            O => \N__35188\,
            I => \current_shift_inst.timer_phase.counter_cry_25\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35185\,
            I => \current_shift_inst.timer_phase.counter_cry_8\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35182\,
            I => \current_shift_inst.timer_phase.counter_cry_9\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35179\,
            I => \current_shift_inst.timer_phase.counter_cry_10\
        );

    \I__7198\ : InMux
    port map (
            O => \N__35176\,
            I => \current_shift_inst.timer_phase.counter_cry_11\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35173\,
            I => \current_shift_inst.timer_phase.counter_cry_12\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35170\,
            I => \current_shift_inst.timer_phase.counter_cry_13\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35167\,
            I => \current_shift_inst.timer_phase.counter_cry_14\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35164\,
            I => \bfn_14_24_0_\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35161\,
            I => \current_shift_inst.timer_phase.counter_cry_16\
        );

    \I__7192\ : InMux
    port map (
            O => \N__35158\,
            I => \bfn_14_22_0_\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35155\,
            I => \current_shift_inst.timer_phase.counter_cry_0\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35152\,
            I => \current_shift_inst.timer_phase.counter_cry_1\
        );

    \I__7189\ : InMux
    port map (
            O => \N__35149\,
            I => \current_shift_inst.timer_phase.counter_cry_2\
        );

    \I__7188\ : InMux
    port map (
            O => \N__35146\,
            I => \current_shift_inst.timer_phase.counter_cry_3\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35143\,
            I => \current_shift_inst.timer_phase.counter_cry_4\
        );

    \I__7186\ : InMux
    port map (
            O => \N__35140\,
            I => \current_shift_inst.timer_phase.counter_cry_5\
        );

    \I__7185\ : InMux
    port map (
            O => \N__35137\,
            I => \current_shift_inst.timer_phase.counter_cry_6\
        );

    \I__7184\ : InMux
    port map (
            O => \N__35134\,
            I => \bfn_14_23_0_\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__35131\,
            I => \N__35127\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35122\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35122\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35122\,
            I => \N__35119\
        );

    \I__7179\ : Span4Mux_v
    port map (
            O => \N__35119\,
            I => \N__35114\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35118\,
            I => \N__35111\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35117\,
            I => \N__35108\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__35114\,
            I => \N__35105\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35111\,
            I => \N__35102\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__35108\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__35105\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__7172\ : Odrv12
    port map (
            O => \N__35102\,
            I => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35095\,
            I => \N__35092\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35092\,
            I => \N__35087\
        );

    \I__7169\ : CascadeMux
    port map (
            O => \N__35091\,
            I => \N__35084\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__35090\,
            I => \N__35081\
        );

    \I__7167\ : Span4Mux_v
    port map (
            O => \N__35087\,
            I => \N__35077\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35074\
        );

    \I__7165\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35069\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35069\
        );

    \I__7163\ : Span4Mux_v
    port map (
            O => \N__35077\,
            I => \N__35066\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__35074\,
            I => \N__35063\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__35069\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__7160\ : Odrv4
    port map (
            O => \N__35066\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__7159\ : Odrv12
    port map (
            O => \N__35063\,
            I => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\
        );

    \I__7158\ : CascadeMux
    port map (
            O => \N__35056\,
            I => \N__35051\
        );

    \I__7157\ : InMux
    port map (
            O => \N__35055\,
            I => \N__35047\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35044\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35039\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35039\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__35047\,
            I => \N__35036\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35044\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35039\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__7150\ : Odrv12
    port map (
            O => \N__35036\,
            I => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\
        );

    \I__7149\ : CascadeMux
    port map (
            O => \N__35029\,
            I => \N__35025\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35028\,
            I => \N__35020\
        );

    \I__7147\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35017\
        );

    \I__7146\ : InMux
    port map (
            O => \N__35024\,
            I => \N__35012\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35023\,
            I => \N__35012\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__35020\,
            I => \N__35009\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__35017\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__35012\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__7141\ : Odrv12
    port map (
            O => \N__35009\,
            I => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\
        );

    \I__7140\ : CascadeMux
    port map (
            O => \N__35002\,
            I => \N__34998\
        );

    \I__7139\ : CascadeMux
    port map (
            O => \N__35001\,
            I => \N__34995\
        );

    \I__7138\ : InMux
    port map (
            O => \N__34998\,
            I => \N__34992\
        );

    \I__7137\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34989\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__34992\,
            I => \N__34986\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__34989\,
            I => \N__34981\
        );

    \I__7134\ : Span4Mux_h
    port map (
            O => \N__34986\,
            I => \N__34978\
        );

    \I__7133\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34975\
        );

    \I__7132\ : InMux
    port map (
            O => \N__34984\,
            I => \N__34972\
        );

    \I__7131\ : Span4Mux_v
    port map (
            O => \N__34981\,
            I => \N__34969\
        );

    \I__7130\ : Odrv4
    port map (
            O => \N__34978\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__34975\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__34972\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__7127\ : Odrv4
    port map (
            O => \N__34969\,
            I => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\
        );

    \I__7126\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34955\
        );

    \I__7125\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34952\
        );

    \I__7124\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34949\
        );

    \I__7123\ : LocalMux
    port map (
            O => \N__34955\,
            I => \N__34946\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__34952\,
            I => \N__34943\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__34949\,
            I => \N__34940\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__34946\,
            I => \N__34937\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__34943\,
            I => \N__34932\
        );

    \I__7118\ : Span4Mux_v
    port map (
            O => \N__34940\,
            I => \N__34932\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__34937\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__34932\,
            I => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\
        );

    \I__7115\ : InMux
    port map (
            O => \N__34927\,
            I => \N__34923\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__34926\,
            I => \N__34920\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__34923\,
            I => \N__34917\
        );

    \I__7112\ : InMux
    port map (
            O => \N__34920\,
            I => \N__34914\
        );

    \I__7111\ : Span4Mux_h
    port map (
            O => \N__34917\,
            I => \N__34908\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__34914\,
            I => \N__34908\
        );

    \I__7109\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34905\
        );

    \I__7108\ : Span4Mux_v
    port map (
            O => \N__34908\,
            I => \N__34902\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__34905\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__34902\,
            I => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\
        );

    \I__7105\ : InMux
    port map (
            O => \N__34897\,
            I => \current_shift_inst.z_cry_30\
        );

    \I__7104\ : InMux
    port map (
            O => \N__34894\,
            I => \N__34890\
        );

    \I__7103\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34887\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__34890\,
            I => \N__34884\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__34887\,
            I => \N__34881\
        );

    \I__7100\ : Span4Mux_h
    port map (
            O => \N__34884\,
            I => \N__34876\
        );

    \I__7099\ : Span4Mux_h
    port map (
            O => \N__34881\,
            I => \N__34876\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__34876\,
            I => \current_shift_inst.z_31\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__34873\,
            I => \N__34870\
        );

    \I__7096\ : InMux
    port map (
            O => \N__34870\,
            I => \N__34867\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__34867\,
            I => \N__34862\
        );

    \I__7094\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34858\
        );

    \I__7093\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34855\
        );

    \I__7092\ : Span4Mux_h
    port map (
            O => \N__34862\,
            I => \N__34852\
        );

    \I__7091\ : InMux
    port map (
            O => \N__34861\,
            I => \N__34849\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__34858\,
            I => \N__34846\
        );

    \I__7089\ : LocalMux
    port map (
            O => \N__34855\,
            I => \N__34843\
        );

    \I__7088\ : Odrv4
    port map (
            O => \N__34852\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__34849\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__7086\ : Odrv12
    port map (
            O => \N__34846\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__7085\ : Odrv12
    port map (
            O => \N__34843\,
            I => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\
        );

    \I__7084\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34830\
        );

    \I__7083\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34826\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__34830\,
            I => \N__34823\
        );

    \I__7081\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34820\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__34826\,
            I => \N__34812\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__34823\,
            I => \N__34812\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34812\
        );

    \I__7077\ : InMux
    port map (
            O => \N__34819\,
            I => \N__34809\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__34812\,
            I => \N__34806\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__34809\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__7074\ : Odrv4
    port map (
            O => \N__34806\,
            I => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\
        );

    \I__7073\ : CascadeMux
    port map (
            O => \N__34801\,
            I => \N__34798\
        );

    \I__7072\ : InMux
    port map (
            O => \N__34798\,
            I => \N__34795\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__34795\,
            I => \N__34791\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__34794\,
            I => \N__34788\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__34791\,
            I => \N__34785\
        );

    \I__7068\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34780\
        );

    \I__7067\ : Span4Mux_v
    port map (
            O => \N__34785\,
            I => \N__34777\
        );

    \I__7066\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34774\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34771\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__34780\,
            I => \N__34768\
        );

    \I__7063\ : Odrv4
    port map (
            O => \N__34777\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34774\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__34771\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__34768\,
            I => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\
        );

    \I__7059\ : CascadeMux
    port map (
            O => \N__34759\,
            I => \N__34756\
        );

    \I__7058\ : InMux
    port map (
            O => \N__34756\,
            I => \N__34750\
        );

    \I__7057\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34750\
        );

    \I__7056\ : LocalMux
    port map (
            O => \N__34750\,
            I => \N__34745\
        );

    \I__7055\ : InMux
    port map (
            O => \N__34749\,
            I => \N__34742\
        );

    \I__7054\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34739\
        );

    \I__7053\ : Span4Mux_h
    port map (
            O => \N__34745\,
            I => \N__34736\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__34742\,
            I => \N__34733\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__34739\,
            I => \N__34730\
        );

    \I__7050\ : Odrv4
    port map (
            O => \N__34736\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__7049\ : Odrv12
    port map (
            O => \N__34733\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__7048\ : Odrv12
    port map (
            O => \N__34730\,
            I => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\
        );

    \I__7047\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34719\
        );

    \I__7046\ : CascadeMux
    port map (
            O => \N__34722\,
            I => \N__34715\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__34719\,
            I => \N__34712\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__34718\,
            I => \N__34709\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34715\,
            I => \N__34705\
        );

    \I__7042\ : Span4Mux_h
    port map (
            O => \N__34712\,
            I => \N__34702\
        );

    \I__7041\ : InMux
    port map (
            O => \N__34709\,
            I => \N__34697\
        );

    \I__7040\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34697\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__34705\,
            I => \N__34694\
        );

    \I__7038\ : Odrv4
    port map (
            O => \N__34702\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__34697\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__7036\ : Odrv12
    port map (
            O => \N__34694\,
            I => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\
        );

    \I__7035\ : CascadeMux
    port map (
            O => \N__34687\,
            I => \N__34682\
        );

    \I__7034\ : CascadeMux
    port map (
            O => \N__34686\,
            I => \N__34679\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34676\
        );

    \I__7032\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34673\
        );

    \I__7031\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34670\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__34676\,
            I => \N__34666\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34663\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__34670\,
            I => \N__34660\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34669\,
            I => \N__34657\
        );

    \I__7026\ : Span4Mux_h
    port map (
            O => \N__34666\,
            I => \N__34654\
        );

    \I__7025\ : Span4Mux_v
    port map (
            O => \N__34663\,
            I => \N__34651\
        );

    \I__7024\ : Odrv12
    port map (
            O => \N__34660\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__34657\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__7022\ : Odrv4
    port map (
            O => \N__34654\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__7021\ : Odrv4
    port map (
            O => \N__34651\,
            I => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\
        );

    \I__7020\ : CascadeMux
    port map (
            O => \N__34642\,
            I => \N__34639\
        );

    \I__7019\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34636\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__34636\,
            I => \N__34632\
        );

    \I__7017\ : CascadeMux
    port map (
            O => \N__34635\,
            I => \N__34629\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__34632\,
            I => \N__34624\
        );

    \I__7015\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34621\
        );

    \I__7014\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34616\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34616\
        );

    \I__7012\ : Span4Mux_h
    port map (
            O => \N__34624\,
            I => \N__34611\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__34621\,
            I => \N__34611\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__34616\,
            I => \N__34608\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__34611\,
            I => \N__34605\
        );

    \I__7008\ : Odrv12
    port map (
            O => \N__34608\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__7007\ : Odrv4
    port map (
            O => \N__34605\,
            I => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\
        );

    \I__7006\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34597\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__34597\,
            I => \N__34591\
        );

    \I__7004\ : InMux
    port map (
            O => \N__34596\,
            I => \N__34586\
        );

    \I__7003\ : InMux
    port map (
            O => \N__34595\,
            I => \N__34586\
        );

    \I__7002\ : CascadeMux
    port map (
            O => \N__34594\,
            I => \N__34583\
        );

    \I__7001\ : Span4Mux_v
    port map (
            O => \N__34591\,
            I => \N__34580\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__34586\,
            I => \N__34577\
        );

    \I__6999\ : InMux
    port map (
            O => \N__34583\,
            I => \N__34574\
        );

    \I__6998\ : Span4Mux_h
    port map (
            O => \N__34580\,
            I => \N__34571\
        );

    \I__6997\ : Span4Mux_h
    port map (
            O => \N__34577\,
            I => \N__34568\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__34574\,
            I => \N__34565\
        );

    \I__6995\ : Odrv4
    port map (
            O => \N__34571\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__34568\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__6993\ : Odrv12
    port map (
            O => \N__34565\,
            I => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\
        );

    \I__6992\ : InMux
    port map (
            O => \N__34558\,
            I => \N__34555\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__34555\,
            I => \N__34551\
        );

    \I__6990\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34546\
        );

    \I__6989\ : Span4Mux_h
    port map (
            O => \N__34551\,
            I => \N__34543\
        );

    \I__6988\ : InMux
    port map (
            O => \N__34550\,
            I => \N__34540\
        );

    \I__6987\ : InMux
    port map (
            O => \N__34549\,
            I => \N__34537\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__34546\,
            I => \N__34534\
        );

    \I__6985\ : Sp12to4
    port map (
            O => \N__34543\,
            I => \N__34529\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__34540\,
            I => \N__34529\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__34537\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__6982\ : Odrv12
    port map (
            O => \N__34534\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__6981\ : Odrv12
    port map (
            O => \N__34529\,
            I => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\
        );

    \I__6980\ : InMux
    port map (
            O => \N__34522\,
            I => \N__34516\
        );

    \I__6979\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34516\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__34516\,
            I => \N__34512\
        );

    \I__6977\ : InMux
    port map (
            O => \N__34515\,
            I => \N__34509\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__34512\,
            I => \N__34506\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__34509\,
            I => \N__34500\
        );

    \I__6974\ : Span4Mux_v
    port map (
            O => \N__34506\,
            I => \N__34500\
        );

    \I__6973\ : InMux
    port map (
            O => \N__34505\,
            I => \N__34497\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__34500\,
            I => \N__34494\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__34497\,
            I => \N__34491\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__34494\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__6969\ : Odrv12
    port map (
            O => \N__34491\,
            I => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\
        );

    \I__6968\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34483\
        );

    \I__6967\ : LocalMux
    port map (
            O => \N__34483\,
            I => \N__34480\
        );

    \I__6966\ : Span4Mux_v
    port map (
            O => \N__34480\,
            I => \N__34475\
        );

    \I__6965\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34472\
        );

    \I__6964\ : CascadeMux
    port map (
            O => \N__34478\,
            I => \N__34469\
        );

    \I__6963\ : Span4Mux_h
    port map (
            O => \N__34475\,
            I => \N__34463\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__34472\,
            I => \N__34463\
        );

    \I__6961\ : InMux
    port map (
            O => \N__34469\,
            I => \N__34460\
        );

    \I__6960\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34457\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__34463\,
            I => \N__34454\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__34460\,
            I => \N__34451\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__34457\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__6956\ : Odrv4
    port map (
            O => \N__34454\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__6955\ : Odrv12
    port map (
            O => \N__34451\,
            I => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__6953\ : InMux
    port map (
            O => \N__34441\,
            I => \N__34434\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34440\,
            I => \N__34434\
        );

    \I__6951\ : InMux
    port map (
            O => \N__34439\,
            I => \N__34431\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34428\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__34431\,
            I => \N__34425\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__34428\,
            I => \N__34422\
        );

    \I__6947\ : Span4Mux_h
    port map (
            O => \N__34425\,
            I => \N__34418\
        );

    \I__6946\ : Span4Mux_h
    port map (
            O => \N__34422\,
            I => \N__34415\
        );

    \I__6945\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34412\
        );

    \I__6944\ : Sp12to4
    port map (
            O => \N__34418\,
            I => \N__34405\
        );

    \I__6943\ : Sp12to4
    port map (
            O => \N__34415\,
            I => \N__34405\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__34412\,
            I => \N__34405\
        );

    \I__6941\ : Odrv12
    port map (
            O => \N__34405\,
            I => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\
        );

    \I__6940\ : CascadeMux
    port map (
            O => \N__34402\,
            I => \N__34397\
        );

    \I__6939\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34394\
        );

    \I__6938\ : InMux
    port map (
            O => \N__34400\,
            I => \N__34390\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34397\,
            I => \N__34387\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34394\,
            I => \N__34384\
        );

    \I__6935\ : CascadeMux
    port map (
            O => \N__34393\,
            I => \N__34381\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__34390\,
            I => \N__34378\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34373\
        );

    \I__6932\ : Span4Mux_v
    port map (
            O => \N__34384\,
            I => \N__34373\
        );

    \I__6931\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34370\
        );

    \I__6930\ : Span4Mux_h
    port map (
            O => \N__34378\,
            I => \N__34363\
        );

    \I__6929\ : Span4Mux_h
    port map (
            O => \N__34373\,
            I => \N__34363\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__34370\,
            I => \N__34363\
        );

    \I__6927\ : Span4Mux_v
    port map (
            O => \N__34363\,
            I => \N__34360\
        );

    \I__6926\ : Odrv4
    port map (
            O => \N__34360\,
            I => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\
        );

    \I__6925\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34352\
        );

    \I__6924\ : CascadeMux
    port map (
            O => \N__34356\,
            I => \N__34349\
        );

    \I__6923\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34346\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__34352\,
            I => \N__34343\
        );

    \I__6921\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34340\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__34346\,
            I => \N__34336\
        );

    \I__6919\ : Span4Mux_v
    port map (
            O => \N__34343\,
            I => \N__34333\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__34340\,
            I => \N__34330\
        );

    \I__6917\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34327\
        );

    \I__6916\ : Span4Mux_v
    port map (
            O => \N__34336\,
            I => \N__34324\
        );

    \I__6915\ : Span4Mux_h
    port map (
            O => \N__34333\,
            I => \N__34319\
        );

    \I__6914\ : Span4Mux_v
    port map (
            O => \N__34330\,
            I => \N__34319\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__34327\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__34324\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__34319\,
            I => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34308\
        );

    \I__6909\ : CascadeMux
    port map (
            O => \N__34311\,
            I => \N__34304\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34300\
        );

    \I__6907\ : InMux
    port map (
            O => \N__34307\,
            I => \N__34297\
        );

    \I__6906\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34294\
        );

    \I__6905\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34291\
        );

    \I__6904\ : Span4Mux_v
    port map (
            O => \N__34300\,
            I => \N__34288\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__34297\,
            I => \N__34285\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__34294\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__34291\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__6900\ : Odrv4
    port map (
            O => \N__34288\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__6899\ : Odrv12
    port map (
            O => \N__34285\,
            I => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34272\
        );

    \I__6897\ : InMux
    port map (
            O => \N__34275\,
            I => \N__34269\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__34272\,
            I => \N__34265\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34269\,
            I => \N__34262\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__34268\,
            I => \N__34259\
        );

    \I__6893\ : Span4Mux_v
    port map (
            O => \N__34265\,
            I => \N__34253\
        );

    \I__6892\ : Span4Mux_v
    port map (
            O => \N__34262\,
            I => \N__34253\
        );

    \I__6891\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34250\
        );

    \I__6890\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34247\
        );

    \I__6889\ : Span4Mux_h
    port map (
            O => \N__34253\,
            I => \N__34244\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__34250\,
            I => \N__34241\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34247\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__34244\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__6885\ : Odrv12
    port map (
            O => \N__34241\,
            I => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34234\,
            I => \N__34229\
        );

    \I__6883\ : CascadeMux
    port map (
            O => \N__34233\,
            I => \N__34226\
        );

    \I__6882\ : InMux
    port map (
            O => \N__34232\,
            I => \N__34223\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__34229\,
            I => \N__34220\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34226\,
            I => \N__34216\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34211\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__34220\,
            I => \N__34211\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34219\,
            I => \N__34208\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34216\,
            I => \N__34205\
        );

    \I__6875\ : Span4Mux_h
    port map (
            O => \N__34211\,
            I => \N__34202\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__34208\,
            I => \N__34199\
        );

    \I__6873\ : Odrv4
    port map (
            O => \N__34205\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__6872\ : Odrv4
    port map (
            O => \N__34202\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__6871\ : Odrv12
    port map (
            O => \N__34199\,
            I => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34192\,
            I => \current_shift_inst.un4_control_input_cry_30\
        );

    \I__6869\ : CascadeMux
    port map (
            O => \N__34189\,
            I => \N__34186\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34186\,
            I => \N__34183\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__34183\,
            I => \N__34180\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__34180\,
            I => \N__34177\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__34177\,
            I => \N__34174\
        );

    \I__6864\ : Odrv4
    port map (
            O => \N__34174\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__34171\,
            I => \N__34168\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34165\,
            I => \N__34162\
        );

    \I__6860\ : Span4Mux_v
    port map (
            O => \N__34162\,
            I => \N__34158\
        );

    \I__6859\ : InMux
    port map (
            O => \N__34161\,
            I => \N__34155\
        );

    \I__6858\ : Span4Mux_h
    port map (
            O => \N__34158\,
            I => \N__34150\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__34155\,
            I => \N__34150\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__34150\,
            I => \N__34147\
        );

    \I__6855\ : Odrv4
    port map (
            O => \N__34147\,
            I => \current_shift_inst.un38_control_input_0\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34144\,
            I => \N__34140\
        );

    \I__6853\ : CascadeMux
    port map (
            O => \N__34143\,
            I => \N__34137\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__34140\,
            I => \N__34133\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34137\,
            I => \N__34130\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34136\,
            I => \N__34127\
        );

    \I__6849\ : Span4Mux_v
    port map (
            O => \N__34133\,
            I => \N__34122\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__34130\,
            I => \N__34122\
        );

    \I__6847\ : LocalMux
    port map (
            O => \N__34127\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__34122\,
            I => \current_shift_inst.elapsed_time_ns_1_fast_31\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__34117\,
            I => \N__34114\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34111\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34111\,
            I => \G_407\
        );

    \I__6842\ : InMux
    port map (
            O => \N__34108\,
            I => \N__34104\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34101\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__34104\,
            I => \N__34096\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34101\,
            I => \N__34096\
        );

    \I__6838\ : Span4Mux_v
    port map (
            O => \N__34096\,
            I => \N__34092\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34089\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__34092\,
            I => \N__34084\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34089\,
            I => \N__34084\
        );

    \I__6834\ : Span4Mux_v
    port map (
            O => \N__34084\,
            I => \N__34081\
        );

    \I__6833\ : Odrv4
    port map (
            O => \N__34081\,
            I => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\
        );

    \I__6832\ : CascadeMux
    port map (
            O => \N__34078\,
            I => \N__34075\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34072\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__34072\,
            I => \G_406\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34066\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34066\,
            I => \N__34062\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34059\
        );

    \I__6826\ : Span4Mux_v
    port map (
            O => \N__34062\,
            I => \N__34053\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__34059\,
            I => \N__34053\
        );

    \I__6824\ : CascadeMux
    port map (
            O => \N__34058\,
            I => \N__34050\
        );

    \I__6823\ : Span4Mux_h
    port map (
            O => \N__34053\,
            I => \N__34047\
        );

    \I__6822\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34044\
        );

    \I__6821\ : Span4Mux_v
    port map (
            O => \N__34047\,
            I => \N__34041\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34038\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__34041\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__6818\ : Odrv12
    port map (
            O => \N__34038\,
            I => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\
        );

    \I__6817\ : InMux
    port map (
            O => \N__34033\,
            I => \N__34029\
        );

    \I__6816\ : CascadeMux
    port map (
            O => \N__34032\,
            I => \N__34026\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34029\,
            I => \N__34023\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34020\
        );

    \I__6813\ : Span4Mux_h
    port map (
            O => \N__34023\,
            I => \N__34017\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__34014\
        );

    \I__6811\ : Span4Mux_v
    port map (
            O => \N__34017\,
            I => \N__34009\
        );

    \I__6810\ : Span4Mux_v
    port map (
            O => \N__34014\,
            I => \N__34009\
        );

    \I__6809\ : Odrv4
    port map (
            O => \N__34009\,
            I => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\
        );

    \I__6808\ : CascadeMux
    port map (
            O => \N__34006\,
            I => \N__34003\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33996\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33996\
        );

    \I__6805\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33993\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__33996\,
            I => \N__33990\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33986\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__33990\,
            I => \N__33983\
        );

    \I__6801\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33980\
        );

    \I__6800\ : Span4Mux_v
    port map (
            O => \N__33986\,
            I => \N__33977\
        );

    \I__6799\ : Span4Mux_h
    port map (
            O => \N__33983\,
            I => \N__33974\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__33980\,
            I => \N__33971\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__33977\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__33974\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__6795\ : Odrv12
    port map (
            O => \N__33971\,
            I => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__33964\,
            I => \N__33961\
        );

    \I__6793\ : InMux
    port map (
            O => \N__33961\,
            I => \N__33957\
        );

    \I__6792\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33954\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__33957\,
            I => \N__33950\
        );

    \I__6790\ : LocalMux
    port map (
            O => \N__33954\,
            I => \N__33947\
        );

    \I__6789\ : InMux
    port map (
            O => \N__33953\,
            I => \N__33944\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__33950\,
            I => \N__33936\
        );

    \I__6787\ : Span4Mux_v
    port map (
            O => \N__33947\,
            I => \N__33936\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__33944\,
            I => \N__33936\
        );

    \I__6785\ : CascadeMux
    port map (
            O => \N__33943\,
            I => \N__33933\
        );

    \I__6784\ : Span4Mux_v
    port map (
            O => \N__33936\,
            I => \N__33930\
        );

    \I__6783\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33927\
        );

    \I__6782\ : Span4Mux_h
    port map (
            O => \N__33930\,
            I => \N__33924\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__33927\,
            I => \N__33921\
        );

    \I__6780\ : Odrv4
    port map (
            O => \N__33924\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__6779\ : Odrv12
    port map (
            O => \N__33921\,
            I => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\
        );

    \I__6778\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33909\
        );

    \I__6777\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33909\
        );

    \I__6776\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33906\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__33909\,
            I => \N__33903\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__33906\,
            I => \N__33898\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__33903\,
            I => \N__33898\
        );

    \I__6772\ : Span4Mux_v
    port map (
            O => \N__33898\,
            I => \N__33894\
        );

    \I__6771\ : InMux
    port map (
            O => \N__33897\,
            I => \N__33891\
        );

    \I__6770\ : Span4Mux_v
    port map (
            O => \N__33894\,
            I => \N__33888\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__33891\,
            I => \N__33885\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__33888\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__6767\ : Odrv12
    port map (
            O => \N__33885\,
            I => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\
        );

    \I__6766\ : InMux
    port map (
            O => \N__33880\,
            I => \current_shift_inst.un4_control_input_cry_21\
        );

    \I__6765\ : InMux
    port map (
            O => \N__33877\,
            I => \current_shift_inst.un4_control_input_cry_22\
        );

    \I__6764\ : InMux
    port map (
            O => \N__33874\,
            I => \current_shift_inst.un4_control_input_cry_23\
        );

    \I__6763\ : InMux
    port map (
            O => \N__33871\,
            I => \bfn_14_17_0_\
        );

    \I__6762\ : InMux
    port map (
            O => \N__33868\,
            I => \current_shift_inst.un4_control_input_cry_25\
        );

    \I__6761\ : InMux
    port map (
            O => \N__33865\,
            I => \current_shift_inst.un4_control_input_cry_26\
        );

    \I__6760\ : InMux
    port map (
            O => \N__33862\,
            I => \current_shift_inst.un4_control_input_cry_27\
        );

    \I__6759\ : InMux
    port map (
            O => \N__33859\,
            I => \current_shift_inst.un4_control_input_cry_28\
        );

    \I__6758\ : InMux
    port map (
            O => \N__33856\,
            I => \current_shift_inst.un4_control_input_cry_29\
        );

    \I__6757\ : InMux
    port map (
            O => \N__33853\,
            I => \current_shift_inst.un4_control_input_cry_12\
        );

    \I__6756\ : InMux
    port map (
            O => \N__33850\,
            I => \current_shift_inst.un4_control_input_cry_13\
        );

    \I__6755\ : InMux
    port map (
            O => \N__33847\,
            I => \current_shift_inst.un4_control_input_cry_14\
        );

    \I__6754\ : InMux
    port map (
            O => \N__33844\,
            I => \current_shift_inst.un4_control_input_cry_15\
        );

    \I__6753\ : InMux
    port map (
            O => \N__33841\,
            I => \bfn_14_16_0_\
        );

    \I__6752\ : InMux
    port map (
            O => \N__33838\,
            I => \current_shift_inst.un4_control_input_cry_17\
        );

    \I__6751\ : InMux
    port map (
            O => \N__33835\,
            I => \current_shift_inst.un4_control_input_cry_18\
        );

    \I__6750\ : InMux
    port map (
            O => \N__33832\,
            I => \current_shift_inst.un4_control_input_cry_19\
        );

    \I__6749\ : InMux
    port map (
            O => \N__33829\,
            I => \current_shift_inst.un4_control_input_cry_20\
        );

    \I__6748\ : InMux
    port map (
            O => \N__33826\,
            I => \current_shift_inst.un4_control_input_cry_3\
        );

    \I__6747\ : InMux
    port map (
            O => \N__33823\,
            I => \current_shift_inst.un4_control_input_cry_4\
        );

    \I__6746\ : InMux
    port map (
            O => \N__33820\,
            I => \current_shift_inst.un4_control_input_cry_5\
        );

    \I__6745\ : InMux
    port map (
            O => \N__33817\,
            I => \current_shift_inst.un4_control_input_cry_6\
        );

    \I__6744\ : InMux
    port map (
            O => \N__33814\,
            I => \current_shift_inst.un4_control_input_cry_7\
        );

    \I__6743\ : InMux
    port map (
            O => \N__33811\,
            I => \bfn_14_15_0_\
        );

    \I__6742\ : InMux
    port map (
            O => \N__33808\,
            I => \current_shift_inst.un4_control_input_cry_9\
        );

    \I__6741\ : InMux
    port map (
            O => \N__33805\,
            I => \current_shift_inst.un4_control_input_cry_10\
        );

    \I__6740\ : InMux
    port map (
            O => \N__33802\,
            I => \current_shift_inst.un4_control_input_cry_11\
        );

    \I__6739\ : InMux
    port map (
            O => \N__33799\,
            I => \bfn_14_13_0_\
        );

    \I__6738\ : InMux
    port map (
            O => \N__33796\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__6737\ : InMux
    port map (
            O => \N__33793\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__6736\ : InMux
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__33787\,
            I => \N__33784\
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__33784\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\
        );

    \I__6733\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33776\
        );

    \I__6732\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33773\
        );

    \I__6731\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33770\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__33776\,
            I => \N__33767\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__33773\,
            I => \N__33761\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__33770\,
            I => \N__33761\
        );

    \I__6727\ : Span4Mux_v
    port map (
            O => \N__33767\,
            I => \N__33758\
        );

    \I__6726\ : InMux
    port map (
            O => \N__33766\,
            I => \N__33755\
        );

    \I__6725\ : Span4Mux_h
    port map (
            O => \N__33761\,
            I => \N__33752\
        );

    \I__6724\ : Span4Mux_h
    port map (
            O => \N__33758\,
            I => \N__33749\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__33755\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6722\ : Odrv4
    port map (
            O => \N__33752\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6721\ : Odrv4
    port map (
            O => \N__33749\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__6720\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33739\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__33739\,
            I => \current_shift_inst.un4_control_input_axb_1\
        );

    \I__6718\ : InMux
    port map (
            O => \N__33736\,
            I => \N__33733\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__33733\,
            I => \current_shift_inst.un4_control_input_axb_2\
        );

    \I__6716\ : InMux
    port map (
            O => \N__33730\,
            I => \current_shift_inst.un4_control_input_cry_1\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33727\,
            I => \N__33724\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__33724\,
            I => \current_shift_inst.un4_control_input_axb_3\
        );

    \I__6713\ : InMux
    port map (
            O => \N__33721\,
            I => \current_shift_inst.un4_control_input_cry_2\
        );

    \I__6712\ : InMux
    port map (
            O => \N__33718\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__6711\ : InMux
    port map (
            O => \N__33715\,
            I => \bfn_14_12_0_\
        );

    \I__6710\ : InMux
    port map (
            O => \N__33712\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33709\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__6708\ : InMux
    port map (
            O => \N__33706\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__6707\ : InMux
    port map (
            O => \N__33703\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33700\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33697\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__6704\ : InMux
    port map (
            O => \N__33694\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__33691\,
            I => \phase_controller_slave.stoper_tr.time_passed11_cascade_\
        );

    \I__6702\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33685\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__33685\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__6700\ : InMux
    port map (
            O => \N__33682\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__6699\ : InMux
    port map (
            O => \N__33679\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__6698\ : InMux
    port map (
            O => \N__33676\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__6697\ : InMux
    port map (
            O => \N__33673\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__6696\ : InMux
    port map (
            O => \N__33670\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__6695\ : InMux
    port map (
            O => \N__33667\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__6694\ : IoInMux
    port map (
            O => \N__33664\,
            I => \N__33661\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__33661\,
            I => \N__33658\
        );

    \I__6692\ : Odrv12
    port map (
            O => \N__33658\,
            I => s2_phy_c
        );

    \I__6691\ : CascadeMux
    port map (
            O => \N__33655\,
            I => \N__33652\
        );

    \I__6690\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33640\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33640\
        );

    \I__6688\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33635\
        );

    \I__6687\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33635\
        );

    \I__6686\ : CascadeMux
    port map (
            O => \N__33648\,
            I => \N__33629\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__33647\,
            I => \N__33623\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__33646\,
            I => \N__33617\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__33645\,
            I => \N__33614\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33640\,
            I => \N__33608\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__33635\,
            I => \N__33608\
        );

    \I__6680\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33605\
        );

    \I__6679\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33599\
        );

    \I__6678\ : InMux
    port map (
            O => \N__33632\,
            I => \N__33596\
        );

    \I__6677\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33593\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33590\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__33627\,
            I => \N__33587\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33575\
        );

    \I__6673\ : InMux
    port map (
            O => \N__33623\,
            I => \N__33575\
        );

    \I__6672\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33575\
        );

    \I__6671\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33575\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33620\,
            I => \N__33575\
        );

    \I__6669\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33567\
        );

    \I__6668\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33567\
        );

    \I__6667\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33567\
        );

    \I__6666\ : Span4Mux_v
    port map (
            O => \N__33608\,
            I => \N__33562\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__33605\,
            I => \N__33562\
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__33604\,
            I => \N__33552\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__33603\,
            I => \N__33549\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__33602\,
            I => \N__33546\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33541\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33534\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__33593\,
            I => \N__33534\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__33590\,
            I => \N__33534\
        );

    \I__6657\ : InMux
    port map (
            O => \N__33587\,
            I => \N__33529\
        );

    \I__6656\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33529\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__33575\,
            I => \N__33526\
        );

    \I__6654\ : InMux
    port map (
            O => \N__33574\,
            I => \N__33523\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__33567\,
            I => \N__33520\
        );

    \I__6652\ : Span4Mux_v
    port map (
            O => \N__33562\,
            I => \N__33517\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33561\,
            I => \N__33510\
        );

    \I__6650\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33510\
        );

    \I__6649\ : InMux
    port map (
            O => \N__33559\,
            I => \N__33510\
        );

    \I__6648\ : InMux
    port map (
            O => \N__33558\,
            I => \N__33501\
        );

    \I__6647\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33501\
        );

    \I__6646\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33501\
        );

    \I__6645\ : InMux
    port map (
            O => \N__33555\,
            I => \N__33501\
        );

    \I__6644\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33490\
        );

    \I__6643\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33490\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33490\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33490\
        );

    \I__6640\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33490\
        );

    \I__6639\ : Span4Mux_h
    port map (
            O => \N__33541\,
            I => \N__33485\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__33534\,
            I => \N__33485\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__33529\,
            I => \N__33480\
        );

    \I__6636\ : Span4Mux_h
    port map (
            O => \N__33526\,
            I => \N__33480\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33473\
        );

    \I__6634\ : Span4Mux_h
    port map (
            O => \N__33520\,
            I => \N__33473\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__33517\,
            I => \N__33473\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__33510\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__33501\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__33490\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__33485\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__33480\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__33473\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__6626\ : InMux
    port map (
            O => \N__33460\,
            I => \N__33457\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__33457\,
            I => \N__33452\
        );

    \I__6624\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33449\
        );

    \I__6623\ : InMux
    port map (
            O => \N__33455\,
            I => \N__33446\
        );

    \I__6622\ : Span4Mux_h
    port map (
            O => \N__33452\,
            I => \N__33438\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__33449\,
            I => \N__33433\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33433\
        );

    \I__6619\ : InMux
    port map (
            O => \N__33445\,
            I => \N__33424\
        );

    \I__6618\ : InMux
    port map (
            O => \N__33444\,
            I => \N__33424\
        );

    \I__6617\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33424\
        );

    \I__6616\ : InMux
    port map (
            O => \N__33442\,
            I => \N__33424\
        );

    \I__6615\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33421\
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__33438\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__6613\ : Odrv12
    port map (
            O => \N__33433\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__33424\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__33421\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__6610\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33408\
        );

    \I__6609\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33403\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33400\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33397\
        );

    \I__6606\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33394\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__33403\,
            I => \N__33388\
        );

    \I__6604\ : Span4Mux_h
    port map (
            O => \N__33400\,
            I => \N__33388\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__33397\,
            I => \N__33385\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__33394\,
            I => \N__33382\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33379\
        );

    \I__6600\ : Odrv4
    port map (
            O => \N__33388\,
            I => measured_delay_hc_12
        );

    \I__6599\ : Odrv12
    port map (
            O => \N__33385\,
            I => measured_delay_hc_12
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__33382\,
            I => measured_delay_hc_12
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__33379\,
            I => measured_delay_hc_12
        );

    \I__6596\ : InMux
    port map (
            O => \N__33370\,
            I => \N__33366\
        );

    \I__6595\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33361\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__33366\,
            I => \N__33357\
        );

    \I__6593\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33354\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33351\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__33361\,
            I => \N__33348\
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__33360\,
            I => \N__33345\
        );

    \I__6589\ : Span4Mux_v
    port map (
            O => \N__33357\,
            I => \N__33342\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__33354\,
            I => \N__33339\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__33351\,
            I => \N__33336\
        );

    \I__6586\ : Span4Mux_v
    port map (
            O => \N__33348\,
            I => \N__33333\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33330\
        );

    \I__6584\ : Span4Mux_h
    port map (
            O => \N__33342\,
            I => \N__33327\
        );

    \I__6583\ : Span4Mux_v
    port map (
            O => \N__33339\,
            I => \N__33324\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__33336\,
            I => \N__33319\
        );

    \I__6581\ : Span4Mux_h
    port map (
            O => \N__33333\,
            I => \N__33319\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__33330\,
            I => measured_delay_hc_14
        );

    \I__6579\ : Odrv4
    port map (
            O => \N__33327\,
            I => measured_delay_hc_14
        );

    \I__6578\ : Odrv4
    port map (
            O => \N__33324\,
            I => measured_delay_hc_14
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__33319\,
            I => measured_delay_hc_14
        );

    \I__6576\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33303\
        );

    \I__6575\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33300\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__33308\,
            I => \N__33297\
        );

    \I__6573\ : InMux
    port map (
            O => \N__33307\,
            I => \N__33294\
        );

    \I__6572\ : CascadeMux
    port map (
            O => \N__33306\,
            I => \N__33291\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33288\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__33300\,
            I => \N__33285\
        );

    \I__6569\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33282\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__33294\,
            I => \N__33279\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33276\
        );

    \I__6566\ : Span4Mux_h
    port map (
            O => \N__33288\,
            I => \N__33273\
        );

    \I__6565\ : Span4Mux_v
    port map (
            O => \N__33285\,
            I => \N__33266\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__33282\,
            I => \N__33266\
        );

    \I__6563\ : Span4Mux_v
    port map (
            O => \N__33279\,
            I => \N__33266\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__33276\,
            I => measured_delay_hc_16
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__33273\,
            I => measured_delay_hc_16
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__33266\,
            I => measured_delay_hc_16
        );

    \I__6559\ : InMux
    port map (
            O => \N__33259\,
            I => \N__33255\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33250\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33246\
        );

    \I__6556\ : InMux
    port map (
            O => \N__33254\,
            I => \N__33243\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33253\,
            I => \N__33240\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__33250\,
            I => \N__33237\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33234\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__33246\,
            I => \N__33231\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33226\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__33240\,
            I => \N__33226\
        );

    \I__6549\ : Span4Mux_v
    port map (
            O => \N__33237\,
            I => \N__33223\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__33234\,
            I => \N__33216\
        );

    \I__6547\ : Span4Mux_h
    port map (
            O => \N__33231\,
            I => \N__33216\
        );

    \I__6546\ : Span4Mux_v
    port map (
            O => \N__33226\,
            I => \N__33216\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__33223\,
            I => measured_delay_hc_17
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__33216\,
            I => measured_delay_hc_17
        );

    \I__6543\ : InMux
    port map (
            O => \N__33211\,
            I => \N__33205\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33201\
        );

    \I__6541\ : CascadeMux
    port map (
            O => \N__33209\,
            I => \N__33198\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33208\,
            I => \N__33195\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__33205\,
            I => \N__33192\
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__33204\,
            I => \N__33189\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__33201\,
            I => \N__33186\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33183\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33178\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__33192\,
            I => \N__33178\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33175\
        );

    \I__6532\ : Span4Mux_h
    port map (
            O => \N__33186\,
            I => \N__33170\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__33183\,
            I => \N__33170\
        );

    \I__6530\ : Odrv4
    port map (
            O => \N__33178\,
            I => measured_delay_hc_18
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__33175\,
            I => measured_delay_hc_18
        );

    \I__6528\ : Odrv4
    port map (
            O => \N__33170\,
            I => measured_delay_hc_18
        );

    \I__6527\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33160\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__33160\,
            I => \N__33156\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33152\
        );

    \I__6524\ : Span4Mux_v
    port map (
            O => \N__33156\,
            I => \N__33149\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33146\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__33152\,
            I => \N__33143\
        );

    \I__6521\ : Span4Mux_h
    port map (
            O => \N__33149\,
            I => \N__33140\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__33146\,
            I => \N__33135\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__33143\,
            I => \N__33135\
        );

    \I__6518\ : Odrv4
    port map (
            O => \N__33140\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__33135\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\
        );

    \I__6516\ : InMux
    port map (
            O => \N__33130\,
            I => \N__33126\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33122\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__33126\,
            I => \N__33119\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33116\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__33122\,
            I => \N__33112\
        );

    \I__6511\ : Span4Mux_h
    port map (
            O => \N__33119\,
            I => \N__33109\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__33116\,
            I => \N__33106\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33103\
        );

    \I__6508\ : Span4Mux_v
    port map (
            O => \N__33112\,
            I => \N__33100\
        );

    \I__6507\ : Span4Mux_v
    port map (
            O => \N__33109\,
            I => \N__33097\
        );

    \I__6506\ : Span4Mux_v
    port map (
            O => \N__33106\,
            I => \N__33094\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__33103\,
            I => \N__33091\
        );

    \I__6504\ : Odrv4
    port map (
            O => \N__33100\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__33097\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__33094\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__6501\ : Odrv4
    port map (
            O => \N__33091\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\
        );

    \I__6500\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__33079\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33072\
        );

    \I__6497\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33069\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33066\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33069\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__33066\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33058\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33058\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__33055\,
            I => \N__33051\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33048\
        );

    \I__6489\ : InMux
    port map (
            O => \N__33051\,
            I => \N__33045\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__33048\,
            I => \N__33042\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__33045\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6486\ : Odrv12
    port map (
            O => \N__33042\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__6485\ : InMux
    port map (
            O => \N__33037\,
            I => \N__33034\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__33034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__33031\,
            I => \N__33027\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33024\
        );

    \I__6481\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33021\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__33018\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33021\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6478\ : Odrv12
    port map (
            O => \N__33018\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33013\,
            I => \N__33010\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__33010\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33007\,
            I => \N__33003\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33006\,
            I => \N__33000\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__33003\,
            I => \N__32997\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33000\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6471\ : Odrv12
    port map (
            O => \N__32997\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__6470\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32989\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__32989\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__6468\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32982\
        );

    \I__6467\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32979\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__32982\,
            I => \N__32976\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__32979\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6464\ : Odrv12
    port map (
            O => \N__32976\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__6463\ : InMux
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__32968\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__6461\ : InMux
    port map (
            O => \N__32965\,
            I => \N__32962\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__32962\,
            I => \N__32958\
        );

    \I__6459\ : InMux
    port map (
            O => \N__32961\,
            I => \N__32955\
        );

    \I__6458\ : Span4Mux_v
    port map (
            O => \N__32958\,
            I => \N__32952\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__32955\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__32952\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__6455\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__32944\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__6453\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32937\
        );

    \I__6452\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32934\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__32937\,
            I => \N__32931\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__32934\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__6449\ : Odrv12
    port map (
            O => \N__32931\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__32926\,
            I => \N__32920\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__32925\,
            I => \N__32917\
        );

    \I__6446\ : InMux
    port map (
            O => \N__32924\,
            I => \N__32914\
        );

    \I__6445\ : CascadeMux
    port map (
            O => \N__32923\,
            I => \N__32910\
        );

    \I__6444\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32889\
        );

    \I__6443\ : InMux
    port map (
            O => \N__32917\,
            I => \N__32889\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__32914\,
            I => \N__32886\
        );

    \I__6441\ : InMux
    port map (
            O => \N__32913\,
            I => \N__32869\
        );

    \I__6440\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32869\
        );

    \I__6439\ : InMux
    port map (
            O => \N__32909\,
            I => \N__32869\
        );

    \I__6438\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32869\
        );

    \I__6437\ : InMux
    port map (
            O => \N__32907\,
            I => \N__32869\
        );

    \I__6436\ : InMux
    port map (
            O => \N__32906\,
            I => \N__32869\
        );

    \I__6435\ : InMux
    port map (
            O => \N__32905\,
            I => \N__32869\
        );

    \I__6434\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32869\
        );

    \I__6433\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32858\
        );

    \I__6432\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32858\
        );

    \I__6431\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32858\
        );

    \I__6430\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32858\
        );

    \I__6429\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32858\
        );

    \I__6428\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32853\
        );

    \I__6427\ : InMux
    port map (
            O => \N__32897\,
            I => \N__32853\
        );

    \I__6426\ : InMux
    port map (
            O => \N__32896\,
            I => \N__32848\
        );

    \I__6425\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32843\
        );

    \I__6424\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32843\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32834\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__32886\,
            I => \N__32834\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__32869\,
            I => \N__32834\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__32858\,
            I => \N__32834\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__32853\,
            I => \N__32831\
        );

    \I__6418\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32828\
        );

    \I__6417\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32825\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32822\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32819\
        );

    \I__6414\ : Span4Mux_v
    port map (
            O => \N__32834\,
            I => \N__32814\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__32831\,
            I => \N__32814\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__32828\,
            I => \N__32811\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__32825\,
            I => \N__32805\
        );

    \I__6410\ : Span12Mux_v
    port map (
            O => \N__32822\,
            I => \N__32805\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__32819\,
            I => \N__32800\
        );

    \I__6408\ : Span4Mux_h
    port map (
            O => \N__32814\,
            I => \N__32800\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__32811\,
            I => \N__32797\
        );

    \I__6406\ : InMux
    port map (
            O => \N__32810\,
            I => \N__32794\
        );

    \I__6405\ : Odrv12
    port map (
            O => \N__32805\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__32800\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__32797\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__32794\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32785\,
            I => \N__32782\
        );

    \I__6400\ : LocalMux
    port map (
            O => \N__32782\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__32779\,
            I => \N__32767\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__32778\,
            I => \N__32764\
        );

    \I__6397\ : CascadeMux
    port map (
            O => \N__32777\,
            I => \N__32761\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__32776\,
            I => \N__32754\
        );

    \I__6395\ : CascadeMux
    port map (
            O => \N__32775\,
            I => \N__32751\
        );

    \I__6394\ : CascadeMux
    port map (
            O => \N__32774\,
            I => \N__32748\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__32773\,
            I => \N__32745\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__32772\,
            I => \N__32741\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__32771\,
            I => \N__32738\
        );

    \I__6390\ : CascadeMux
    port map (
            O => \N__32770\,
            I => \N__32734\
        );

    \I__6389\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32718\
        );

    \I__6388\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32718\
        );

    \I__6387\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32718\
        );

    \I__6386\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32718\
        );

    \I__6385\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32718\
        );

    \I__6384\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32718\
        );

    \I__6383\ : InMux
    port map (
            O => \N__32757\,
            I => \N__32715\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32754\,
            I => \N__32712\
        );

    \I__6381\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32703\
        );

    \I__6380\ : InMux
    port map (
            O => \N__32748\,
            I => \N__32703\
        );

    \I__6379\ : InMux
    port map (
            O => \N__32745\,
            I => \N__32703\
        );

    \I__6378\ : InMux
    port map (
            O => \N__32744\,
            I => \N__32703\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32694\
        );

    \I__6376\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32694\
        );

    \I__6375\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32694\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32734\,
            I => \N__32694\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__32733\,
            I => \N__32691\
        );

    \I__6372\ : CascadeMux
    port map (
            O => \N__32732\,
            I => \N__32687\
        );

    \I__6371\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32681\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__32718\,
            I => \N__32678\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__32715\,
            I => \N__32669\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32669\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32669\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__32694\,
            I => \N__32669\
        );

    \I__6365\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32666\
        );

    \I__6364\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32661\
        );

    \I__6363\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32661\
        );

    \I__6362\ : InMux
    port map (
            O => \N__32686\,
            I => \N__32656\
        );

    \I__6361\ : InMux
    port map (
            O => \N__32685\,
            I => \N__32656\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__32684\,
            I => \N__32653\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32650\
        );

    \I__6358\ : Span4Mux_v
    port map (
            O => \N__32678\,
            I => \N__32645\
        );

    \I__6357\ : Span4Mux_v
    port map (
            O => \N__32669\,
            I => \N__32645\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__32666\,
            I => \N__32642\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32639\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32656\,
            I => \N__32636\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32633\
        );

    \I__6352\ : Span4Mux_v
    port map (
            O => \N__32650\,
            I => \N__32630\
        );

    \I__6351\ : Span4Mux_v
    port map (
            O => \N__32645\,
            I => \N__32627\
        );

    \I__6350\ : Span4Mux_h
    port map (
            O => \N__32642\,
            I => \N__32623\
        );

    \I__6349\ : Span4Mux_v
    port map (
            O => \N__32639\,
            I => \N__32620\
        );

    \I__6348\ : Span12Mux_v
    port map (
            O => \N__32636\,
            I => \N__32617\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__32633\,
            I => \N__32610\
        );

    \I__6346\ : Span4Mux_v
    port map (
            O => \N__32630\,
            I => \N__32610\
        );

    \I__6345\ : Span4Mux_v
    port map (
            O => \N__32627\,
            I => \N__32610\
        );

    \I__6344\ : InMux
    port map (
            O => \N__32626\,
            I => \N__32607\
        );

    \I__6343\ : Odrv4
    port map (
            O => \N__32623\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__32620\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6341\ : Odrv12
    port map (
            O => \N__32617\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6340\ : Odrv4
    port map (
            O => \N__32610\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__32607\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__32596\,
            I => \N__32591\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__32595\,
            I => \N__32587\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__32594\,
            I => \N__32577\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32565\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32548\
        );

    \I__6333\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32548\
        );

    \I__6332\ : InMux
    port map (
            O => \N__32586\,
            I => \N__32548\
        );

    \I__6331\ : InMux
    port map (
            O => \N__32585\,
            I => \N__32548\
        );

    \I__6330\ : InMux
    port map (
            O => \N__32584\,
            I => \N__32548\
        );

    \I__6329\ : InMux
    port map (
            O => \N__32583\,
            I => \N__32548\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32548\
        );

    \I__6327\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32548\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32545\
        );

    \I__6325\ : InMux
    port map (
            O => \N__32577\,
            I => \N__32530\
        );

    \I__6324\ : InMux
    port map (
            O => \N__32576\,
            I => \N__32530\
        );

    \I__6323\ : InMux
    port map (
            O => \N__32575\,
            I => \N__32530\
        );

    \I__6322\ : InMux
    port map (
            O => \N__32574\,
            I => \N__32530\
        );

    \I__6321\ : InMux
    port map (
            O => \N__32573\,
            I => \N__32530\
        );

    \I__6320\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32530\
        );

    \I__6319\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32530\
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__32570\,
            I => \N__32527\
        );

    \I__6317\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32521\
        );

    \I__6316\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32521\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__32565\,
            I => \N__32518\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__32548\,
            I => \N__32515\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32510\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__32530\,
            I => \N__32510\
        );

    \I__6311\ : InMux
    port map (
            O => \N__32527\,
            I => \N__32506\
        );

    \I__6310\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32503\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__32521\,
            I => \N__32500\
        );

    \I__6308\ : Span4Mux_v
    port map (
            O => \N__32518\,
            I => \N__32492\
        );

    \I__6307\ : Span4Mux_v
    port map (
            O => \N__32515\,
            I => \N__32492\
        );

    \I__6306\ : Span4Mux_v
    port map (
            O => \N__32510\,
            I => \N__32492\
        );

    \I__6305\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32489\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__32506\,
            I => \N__32484\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__32503\,
            I => \N__32484\
        );

    \I__6302\ : Span4Mux_h
    port map (
            O => \N__32500\,
            I => \N__32481\
        );

    \I__6301\ : InMux
    port map (
            O => \N__32499\,
            I => \N__32478\
        );

    \I__6300\ : Span4Mux_h
    port map (
            O => \N__32492\,
            I => \N__32473\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__32489\,
            I => \N__32473\
        );

    \I__6298\ : Span4Mux_v
    port map (
            O => \N__32484\,
            I => \N__32469\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__32481\,
            I => \N__32466\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__32478\,
            I => \N__32461\
        );

    \I__6295\ : Span4Mux_v
    port map (
            O => \N__32473\,
            I => \N__32461\
        );

    \I__6294\ : InMux
    port map (
            O => \N__32472\,
            I => \N__32458\
        );

    \I__6293\ : Span4Mux_h
    port map (
            O => \N__32469\,
            I => \N__32453\
        );

    \I__6292\ : Span4Mux_v
    port map (
            O => \N__32466\,
            I => \N__32453\
        );

    \I__6291\ : Span4Mux_v
    port map (
            O => \N__32461\,
            I => \N__32450\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__32458\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__32453\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__6288\ : Odrv4
    port map (
            O => \N__32450\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32443\,
            I => \N__32439\
        );

    \I__6286\ : InMux
    port map (
            O => \N__32442\,
            I => \N__32436\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__32439\,
            I => \N__32433\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__32436\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6283\ : Odrv4
    port map (
            O => \N__32433\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6282\ : InMux
    port map (
            O => \N__32428\,
            I => \N__32425\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__32425\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__6280\ : InMux
    port map (
            O => \N__32422\,
            I => \N__32418\
        );

    \I__6279\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32415\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32412\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__32415\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__32412\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__6275\ : InMux
    port map (
            O => \N__32407\,
            I => \N__32403\
        );

    \I__6274\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32398\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__32403\,
            I => \N__32395\
        );

    \I__6272\ : InMux
    port map (
            O => \N__32402\,
            I => \N__32392\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32401\,
            I => \N__32389\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__32398\,
            I => \N__32386\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__32395\,
            I => \N__32379\
        );

    \I__6268\ : LocalMux
    port map (
            O => \N__32392\,
            I => \N__32379\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__32389\,
            I => \N__32379\
        );

    \I__6266\ : Span4Mux_h
    port map (
            O => \N__32386\,
            I => \N__32376\
        );

    \I__6265\ : Span4Mux_h
    port map (
            O => \N__32379\,
            I => \N__32373\
        );

    \I__6264\ : Odrv4
    port map (
            O => \N__32376\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__6263\ : Odrv4
    port map (
            O => \N__32373\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__6262\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32364\
        );

    \I__6261\ : InMux
    port map (
            O => \N__32367\,
            I => \N__32361\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__32364\,
            I => \N__32357\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32354\
        );

    \I__6258\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32351\
        );

    \I__6257\ : Span4Mux_v
    port map (
            O => \N__32357\,
            I => \N__32345\
        );

    \I__6256\ : Span12Mux_h
    port map (
            O => \N__32354\,
            I => \N__32342\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32339\
        );

    \I__6254\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32336\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32349\,
            I => \N__32331\
        );

    \I__6252\ : InMux
    port map (
            O => \N__32348\,
            I => \N__32331\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__32345\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6250\ : Odrv12
    port map (
            O => \N__32342\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6249\ : Odrv12
    port map (
            O => \N__32339\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__32336\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__32331\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__6246\ : CascadeMux
    port map (
            O => \N__32320\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\
        );

    \I__6245\ : CascadeMux
    port map (
            O => \N__32317\,
            I => \N__32312\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32316\,
            I => \N__32309\
        );

    \I__6243\ : InMux
    port map (
            O => \N__32315\,
            I => \N__32306\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32303\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__32309\,
            I => \N__32300\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__32306\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__32303\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6238\ : Odrv4
    port map (
            O => \N__32300\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6237\ : InMux
    port map (
            O => \N__32293\,
            I => \N__32290\
        );

    \I__6236\ : LocalMux
    port map (
            O => \N__32290\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__6235\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32283\
        );

    \I__6234\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32280\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__32283\,
            I => \N__32277\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__32280\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__6231\ : Odrv4
    port map (
            O => \N__32277\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__6230\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32269\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__32269\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32266\,
            I => \N__32262\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32265\,
            I => \N__32259\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32256\
        );

    \I__6225\ : LocalMux
    port map (
            O => \N__32259\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__32256\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__6223\ : InMux
    port map (
            O => \N__32251\,
            I => \N__32248\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__32248\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32245\,
            I => \N__32241\
        );

    \I__6220\ : InMux
    port map (
            O => \N__32244\,
            I => \N__32238\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__32241\,
            I => \N__32235\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__32238\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__6217\ : Odrv4
    port map (
            O => \N__32235\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__6216\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32227\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32227\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__6214\ : InMux
    port map (
            O => \N__32224\,
            I => \N__32220\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32217\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__32220\,
            I => \N__32214\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__32217\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__32214\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32206\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32206\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32199\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32202\,
            I => \N__32196\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__32199\,
            I => \N__32193\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__32196\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__6203\ : Odrv4
    port map (
            O => \N__32193\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32188\,
            I => \N__32185\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__32185\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__6200\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32178\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32175\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__32178\,
            I => \N__32172\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__32175\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__32172\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__6195\ : CascadeMux
    port map (
            O => \N__32167\,
            I => \N__32164\
        );

    \I__6194\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32161\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32161\,
            I => \N__32158\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__32158\,
            I => \N__32155\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__32155\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__6190\ : InMux
    port map (
            O => \N__32152\,
            I => \N__32149\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32149\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__6188\ : InMux
    port map (
            O => \N__32146\,
            I => \N__32142\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__32145\,
            I => \N__32139\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32142\,
            I => \N__32136\
        );

    \I__6185\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32133\
        );

    \I__6184\ : Span4Mux_h
    port map (
            O => \N__32136\,
            I => \N__32130\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__32133\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__32130\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6181\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32122\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32122\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__6179\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32116\
        );

    \I__6178\ : LocalMux
    port map (
            O => \N__32116\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__32113\,
            I => \N__32110\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32107\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32107\,
            I => \N__32104\
        );

    \I__6174\ : Odrv12
    port map (
            O => \N__32104\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32098\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__32098\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__6171\ : InMux
    port map (
            O => \N__32095\,
            I => \N__32092\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__32092\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__6169\ : InMux
    port map (
            O => \N__32089\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__32086\,
            I => \N__32083\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32080\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__32080\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__6165\ : CascadeMux
    port map (
            O => \N__32077\,
            I => \N__32074\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32071\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32071\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__32068\,
            I => \N__32065\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32065\,
            I => \N__32062\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__32062\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__6159\ : InMux
    port map (
            O => \N__32059\,
            I => \N__32056\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__32056\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__6157\ : CascadeMux
    port map (
            O => \N__32053\,
            I => \N__32050\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32047\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32047\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__6154\ : InMux
    port map (
            O => \N__32044\,
            I => \N__32040\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32043\,
            I => \N__32037\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32040\,
            I => \N__32034\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32031\
        );

    \I__6150\ : Odrv12
    port map (
            O => \N__32034\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__32031\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32026\,
            I => \N__32023\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__32023\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__32020\,
            I => \N__32017\
        );

    \I__6145\ : InMux
    port map (
            O => \N__32017\,
            I => \N__32014\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32014\,
            I => \N__32011\
        );

    \I__6143\ : Odrv4
    port map (
            O => \N__32011\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32008\,
            I => \N__32004\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32001\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__31998\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31995\
        );

    \I__6138\ : Odrv12
    port map (
            O => \N__31998\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__6137\ : Odrv4
    port map (
            O => \N__31995\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__6136\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31987\
        );

    \I__6135\ : LocalMux
    port map (
            O => \N__31987\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__6134\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31981\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__31981\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__6132\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31975\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__31975\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__6130\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31969\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__31969\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__6128\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31963\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__31963\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__6126\ : CascadeMux
    port map (
            O => \N__31960\,
            I => \N__31957\
        );

    \I__6125\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31954\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31951\
        );

    \I__6123\ : Odrv4
    port map (
            O => \N__31951\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__6122\ : InMux
    port map (
            O => \N__31948\,
            I => \N__31945\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__31945\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__6120\ : CascadeMux
    port map (
            O => \N__31942\,
            I => \N__31939\
        );

    \I__6119\ : InMux
    port map (
            O => \N__31939\,
            I => \N__31936\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31933\
        );

    \I__6117\ : Span4Mux_v
    port map (
            O => \N__31933\,
            I => \N__31930\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__31930\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__6115\ : InMux
    port map (
            O => \N__31927\,
            I => \N__31924\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__31924\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__31921\,
            I => \N__31918\
        );

    \I__6112\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31915\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__31915\,
            I => \N__31912\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__31912\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__6109\ : InMux
    port map (
            O => \N__31909\,
            I => \N__31906\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__31906\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__6107\ : CascadeMux
    port map (
            O => \N__31903\,
            I => \N__31900\
        );

    \I__6106\ : InMux
    port map (
            O => \N__31900\,
            I => \N__31897\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__31897\,
            I => \N__31894\
        );

    \I__6104\ : Odrv12
    port map (
            O => \N__31894\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__6103\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31888\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__31888\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__6101\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31882\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__31882\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__31879\,
            I => \N__31876\
        );

    \I__6098\ : InMux
    port map (
            O => \N__31876\,
            I => \N__31873\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__31873\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__6096\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31867\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__31867\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__31864\,
            I => \N__31861\
        );

    \I__6093\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31858\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__31858\,
            I => \N__31855\
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__31855\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__6090\ : InMux
    port map (
            O => \N__31852\,
            I => \N__31849\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__31849\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__6088\ : InMux
    port map (
            O => \N__31846\,
            I => \N__31841\
        );

    \I__6087\ : InMux
    port map (
            O => \N__31845\,
            I => \N__31838\
        );

    \I__6086\ : InMux
    port map (
            O => \N__31844\,
            I => \N__31835\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__31841\,
            I => \N__31832\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__31838\,
            I => \N__31826\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31826\
        );

    \I__6082\ : Span4Mux_h
    port map (
            O => \N__31832\,
            I => \N__31823\
        );

    \I__6081\ : InMux
    port map (
            O => \N__31831\,
            I => \N__31820\
        );

    \I__6080\ : Span4Mux_v
    port map (
            O => \N__31826\,
            I => \N__31817\
        );

    \I__6079\ : Span4Mux_v
    port map (
            O => \N__31823\,
            I => \N__31814\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__31820\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6077\ : Odrv4
    port map (
            O => \N__31817\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6076\ : Odrv4
    port map (
            O => \N__31814\,
            I => \current_shift_inst.timer_phase.runningZ0\
        );

    \I__6075\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31804\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31801\
        );

    \I__6073\ : Span4Mux_h
    port map (
            O => \N__31801\,
            I => \N__31798\
        );

    \I__6072\ : Span4Mux_v
    port map (
            O => \N__31798\,
            I => \N__31795\
        );

    \I__6071\ : Odrv4
    port map (
            O => \N__31795\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\
        );

    \I__6070\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31788\
        );

    \I__6069\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31785\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__31788\,
            I => \N__31781\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__31785\,
            I => \N__31778\
        );

    \I__6066\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31775\
        );

    \I__6065\ : Span4Mux_v
    port map (
            O => \N__31781\,
            I => \N__31772\
        );

    \I__6064\ : Span4Mux_v
    port map (
            O => \N__31778\,
            I => \N__31769\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__31775\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6062\ : Odrv4
    port map (
            O => \N__31772\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6061\ : Odrv4
    port map (
            O => \N__31769\,
            I => \current_shift_inst.start_timer_phaseZ0\
        );

    \I__6060\ : InMux
    port map (
            O => \N__31762\,
            I => \N__31757\
        );

    \I__6059\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31754\
        );

    \I__6058\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31751\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__31757\,
            I => \N__31747\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31744\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__31751\,
            I => \N__31741\
        );

    \I__6054\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31738\
        );

    \I__6053\ : Span12Mux_h
    port map (
            O => \N__31747\,
            I => \N__31735\
        );

    \I__6052\ : Span12Mux_v
    port map (
            O => \N__31744\,
            I => \N__31732\
        );

    \I__6051\ : Span4Mux_h
    port map (
            O => \N__31741\,
            I => \N__31729\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__31738\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6049\ : Odrv12
    port map (
            O => \N__31735\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6048\ : Odrv12
    port map (
            O => \N__31732\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__31729\,
            I => \current_shift_inst.stop_timer_phaseZ0\
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__31720\,
            I => \N__31717\
        );

    \I__6045\ : InMux
    port map (
            O => \N__31717\,
            I => \N__31714\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__31714\,
            I => \N__31711\
        );

    \I__6043\ : Span4Mux_v
    port map (
            O => \N__31711\,
            I => \N__31708\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__31708\,
            I => \N__31705\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__31705\,
            I => \N__31702\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__31702\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__31699\,
            I => \N__31696\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31696\,
            I => \N__31693\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__31693\,
            I => \N__31690\
        );

    \I__6036\ : Span4Mux_v
    port map (
            O => \N__31690\,
            I => \N__31687\
        );

    \I__6035\ : Span4Mux_v
    port map (
            O => \N__31687\,
            I => \N__31684\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__31684\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\
        );

    \I__6033\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31678\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__31678\,
            I => \N__31675\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__31675\,
            I => \N__31672\
        );

    \I__6030\ : Span4Mux_v
    port map (
            O => \N__31672\,
            I => \N__31669\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__31669\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\
        );

    \I__6028\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31663\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__31663\,
            I => \N__31660\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__31660\,
            I => \N__31657\
        );

    \I__6025\ : Span4Mux_v
    port map (
            O => \N__31657\,
            I => \N__31654\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__31654\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\
        );

    \I__6023\ : InMux
    port map (
            O => \N__31651\,
            I => \N__31648\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__31648\,
            I => \N__31645\
        );

    \I__6021\ : Span4Mux_v
    port map (
            O => \N__31645\,
            I => \N__31642\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__31642\,
            I => \N__31639\
        );

    \I__6019\ : Odrv4
    port map (
            O => \N__31639\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\
        );

    \I__6018\ : InMux
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__31633\,
            I => \N__31630\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__31630\,
            I => \N__31627\
        );

    \I__6015\ : Span4Mux_v
    port map (
            O => \N__31627\,
            I => \N__31624\
        );

    \I__6014\ : Odrv4
    port map (
            O => \N__31624\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\
        );

    \I__6013\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31618\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__31618\,
            I => \N__31615\
        );

    \I__6011\ : Span4Mux_v
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__31612\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\
        );

    \I__6009\ : CascadeMux
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__6008\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__6005\ : Span4Mux_h
    port map (
            O => \N__31597\,
            I => \N__31594\
        );

    \I__6004\ : Span4Mux_v
    port map (
            O => \N__31594\,
            I => \N__31591\
        );

    \I__6003\ : Odrv4
    port map (
            O => \N__31591\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\
        );

    \I__6002\ : InMux
    port map (
            O => \N__31588\,
            I => \N__31585\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__31585\,
            I => \N__31582\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__5999\ : Span4Mux_v
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__31576\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__31573\,
            I => \N__31570\
        );

    \I__5996\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31567\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31567\,
            I => \N__31564\
        );

    \I__5994\ : Span4Mux_v
    port map (
            O => \N__31564\,
            I => \N__31561\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__31561\,
            I => \N__31558\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__31558\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\
        );

    \I__5991\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31552\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__31552\,
            I => \N__31549\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__31549\,
            I => \N__31546\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__31546\,
            I => \N__31543\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__31543\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\
        );

    \I__5986\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31537\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__31537\,
            I => \N__31534\
        );

    \I__5984\ : Span4Mux_h
    port map (
            O => \N__31534\,
            I => \N__31531\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__31531\,
            I => \N__31528\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__31528\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\
        );

    \I__5981\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31522\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__31522\,
            I => \N__31519\
        );

    \I__5979\ : Span4Mux_h
    port map (
            O => \N__31519\,
            I => \N__31516\
        );

    \I__5978\ : Span4Mux_v
    port map (
            O => \N__31516\,
            I => \N__31513\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__31513\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\
        );

    \I__5976\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31507\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__31507\,
            I => \N__31504\
        );

    \I__5974\ : Span4Mux_h
    port map (
            O => \N__31504\,
            I => \N__31501\
        );

    \I__5973\ : Span4Mux_v
    port map (
            O => \N__31501\,
            I => \N__31498\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__31498\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31495\,
            I => \N__31492\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__31492\,
            I => \N__31489\
        );

    \I__5969\ : Span12Mux_h
    port map (
            O => \N__31489\,
            I => \N__31486\
        );

    \I__5968\ : Odrv12
    port map (
            O => \N__31486\,
            I => \current_shift_inst.un38_control_input_0_axb_31\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__31483\,
            I => \N__31480\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31480\,
            I => \N__31477\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__31477\,
            I => \N__31474\
        );

    \I__5964\ : Span4Mux_h
    port map (
            O => \N__31474\,
            I => \N__31471\
        );

    \I__5963\ : Span4Mux_v
    port map (
            O => \N__31471\,
            I => \N__31468\
        );

    \I__5962\ : Odrv4
    port map (
            O => \N__31468\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\
        );

    \I__5961\ : CEMux
    port map (
            O => \N__31465\,
            I => \N__31461\
        );

    \I__5960\ : CEMux
    port map (
            O => \N__31464\,
            I => \N__31458\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__31461\,
            I => \N__31455\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__31458\,
            I => \N__31451\
        );

    \I__5957\ : Span4Mux_v
    port map (
            O => \N__31455\,
            I => \N__31448\
        );

    \I__5956\ : CEMux
    port map (
            O => \N__31454\,
            I => \N__31445\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__31451\,
            I => \N__31441\
        );

    \I__5954\ : Span4Mux_v
    port map (
            O => \N__31448\,
            I => \N__31436\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31436\
        );

    \I__5952\ : CEMux
    port map (
            O => \N__31444\,
            I => \N__31433\
        );

    \I__5951\ : Span4Mux_h
    port map (
            O => \N__31441\,
            I => \N__31424\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__31436\,
            I => \N__31424\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__31433\,
            I => \N__31424\
        );

    \I__5948\ : CEMux
    port map (
            O => \N__31432\,
            I => \N__31421\
        );

    \I__5947\ : IoInMux
    port map (
            O => \N__31431\,
            I => \N__31418\
        );

    \I__5946\ : Span4Mux_v
    port map (
            O => \N__31424\,
            I => \N__31413\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__31421\,
            I => \N__31413\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__31418\,
            I => \N__31409\
        );

    \I__5943\ : Span4Mux_v
    port map (
            O => \N__31413\,
            I => \N__31406\
        );

    \I__5942\ : CEMux
    port map (
            O => \N__31412\,
            I => \N__31403\
        );

    \I__5941\ : Span4Mux_s1_v
    port map (
            O => \N__31409\,
            I => \N__31400\
        );

    \I__5940\ : Sp12to4
    port map (
            O => \N__31406\,
            I => \N__31395\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__31403\,
            I => \N__31395\
        );

    \I__5938\ : Span4Mux_h
    port map (
            O => \N__31400\,
            I => \N__31392\
        );

    \I__5937\ : Odrv12
    port map (
            O => \N__31395\,
            I => red_c_i
        );

    \I__5936\ : Odrv4
    port map (
            O => \N__31392\,
            I => red_c_i
        );

    \I__5935\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31384\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__31384\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\
        );

    \I__5933\ : InMux
    port map (
            O => \N__31381\,
            I => \N__31378\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__31378\,
            I => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\
        );

    \I__5931\ : CascadeMux
    port map (
            O => \N__31375\,
            I => \N__31372\
        );

    \I__5930\ : InMux
    port map (
            O => \N__31372\,
            I => \N__31369\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__31369\,
            I => \N__31366\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__31366\,
            I => \N__31363\
        );

    \I__5927\ : Span4Mux_v
    port map (
            O => \N__31363\,
            I => \N__31360\
        );

    \I__5926\ : Odrv4
    port map (
            O => \N__31360\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__31357\,
            I => \N__31352\
        );

    \I__5924\ : CascadeMux
    port map (
            O => \N__31356\,
            I => \N__31349\
        );

    \I__5923\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31346\
        );

    \I__5922\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31341\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31341\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__31346\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__31341\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__5918\ : InMux
    port map (
            O => \N__31336\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__5917\ : InMux
    port map (
            O => \N__31333\,
            I => \N__31328\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31332\,
            I => \N__31325\
        );

    \I__5915\ : InMux
    port map (
            O => \N__31331\,
            I => \N__31322\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__31328\,
            I => \N__31319\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__31325\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__31322\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__31319\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__5910\ : InMux
    port map (
            O => \N__31312\,
            I => \bfn_13_10_0_\
        );

    \I__5909\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31304\
        );

    \I__5908\ : InMux
    port map (
            O => \N__31308\,
            I => \N__31301\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31298\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__31304\,
            I => \N__31295\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__31301\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__31298\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__31295\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__5902\ : InMux
    port map (
            O => \N__31288\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__31285\,
            I => \N__31280\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__31284\,
            I => \N__31277\
        );

    \I__5899\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31274\
        );

    \I__5898\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31269\
        );

    \I__5897\ : InMux
    port map (
            O => \N__31277\,
            I => \N__31269\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__31274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__31269\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31264\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__31261\,
            I => \N__31256\
        );

    \I__5892\ : CascadeMux
    port map (
            O => \N__31260\,
            I => \N__31253\
        );

    \I__5891\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31250\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31245\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31253\,
            I => \N__31245\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__31250\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__31245\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__5886\ : InMux
    port map (
            O => \N__31240\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__5885\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31233\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31230\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31233\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__31230\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31225\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__5880\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31188\
        );

    \I__5879\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31188\
        );

    \I__5878\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31179\
        );

    \I__5877\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31179\
        );

    \I__5876\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31179\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31179\
        );

    \I__5874\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31170\
        );

    \I__5873\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31170\
        );

    \I__5872\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31170\
        );

    \I__5871\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31170\
        );

    \I__5870\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31161\
        );

    \I__5869\ : InMux
    port map (
            O => \N__31211\,
            I => \N__31161\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31210\,
            I => \N__31161\
        );

    \I__5867\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31161\
        );

    \I__5866\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31152\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31207\,
            I => \N__31152\
        );

    \I__5864\ : InMux
    port map (
            O => \N__31206\,
            I => \N__31152\
        );

    \I__5863\ : InMux
    port map (
            O => \N__31205\,
            I => \N__31152\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31204\,
            I => \N__31143\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31203\,
            I => \N__31143\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31143\
        );

    \I__5859\ : InMux
    port map (
            O => \N__31201\,
            I => \N__31143\
        );

    \I__5858\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31134\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31199\,
            I => \N__31134\
        );

    \I__5856\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31134\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31134\
        );

    \I__5854\ : InMux
    port map (
            O => \N__31196\,
            I => \N__31125\
        );

    \I__5853\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31125\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31125\
        );

    \I__5851\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31125\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__31188\,
            I => \N__31116\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31116\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__31170\,
            I => \N__31116\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__31161\,
            I => \N__31116\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__31152\,
            I => \N__31109\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31143\,
            I => \N__31109\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31134\,
            I => \N__31109\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__31125\,
            I => \N__31104\
        );

    \I__5842\ : Span4Mux_v
    port map (
            O => \N__31116\,
            I => \N__31104\
        );

    \I__5841\ : Odrv12
    port map (
            O => \N__31109\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__31104\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__5839\ : InMux
    port map (
            O => \N__31099\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__5838\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31092\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__31092\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__31089\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__5834\ : CEMux
    port map (
            O => \N__31084\,
            I => \N__31079\
        );

    \I__5833\ : CEMux
    port map (
            O => \N__31083\,
            I => \N__31076\
        );

    \I__5832\ : CEMux
    port map (
            O => \N__31082\,
            I => \N__31073\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__31079\,
            I => \N__31069\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31076\,
            I => \N__31066\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31063\
        );

    \I__5828\ : CEMux
    port map (
            O => \N__31072\,
            I => \N__31060\
        );

    \I__5827\ : Span4Mux_v
    port map (
            O => \N__31069\,
            I => \N__31055\
        );

    \I__5826\ : Span4Mux_h
    port map (
            O => \N__31066\,
            I => \N__31055\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__31063\,
            I => \N__31052\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__31049\
        );

    \I__5823\ : Span4Mux_h
    port map (
            O => \N__31055\,
            I => \N__31046\
        );

    \I__5822\ : Span4Mux_h
    port map (
            O => \N__31052\,
            I => \N__31043\
        );

    \I__5821\ : Span4Mux_h
    port map (
            O => \N__31049\,
            I => \N__31040\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__31046\,
            I => \delay_measurement_inst.delay_hc_timer.N_337_i\
        );

    \I__5819\ : Odrv4
    port map (
            O => \N__31043\,
            I => \delay_measurement_inst.delay_hc_timer.N_337_i\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__31040\,
            I => \delay_measurement_inst.delay_hc_timer.N_337_i\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__31033\,
            I => \N__31029\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31032\,
            I => \N__31025\
        );

    \I__5815\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31022\
        );

    \I__5814\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31018\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__31025\,
            I => \N__31015\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__31022\,
            I => \N__31012\
        );

    \I__5811\ : InMux
    port map (
            O => \N__31021\,
            I => \N__31009\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__31018\,
            I => \N__31005\
        );

    \I__5809\ : Span4Mux_v
    port map (
            O => \N__31015\,
            I => \N__31002\
        );

    \I__5808\ : Span4Mux_h
    port map (
            O => \N__31012\,
            I => \N__30999\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__31009\,
            I => \N__30996\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31008\,
            I => \N__30993\
        );

    \I__5805\ : Span4Mux_s3_v
    port map (
            O => \N__31005\,
            I => \N__30989\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__31002\,
            I => \N__30985\
        );

    \I__5803\ : Span4Mux_h
    port map (
            O => \N__30999\,
            I => \N__30977\
        );

    \I__5802\ : Span4Mux_v
    port map (
            O => \N__30996\,
            I => \N__30977\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30977\
        );

    \I__5800\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30974\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__30989\,
            I => \N__30971\
        );

    \I__5798\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30968\
        );

    \I__5797\ : Sp12to4
    port map (
            O => \N__30985\,
            I => \N__30965\
        );

    \I__5796\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30962\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__30977\,
            I => \N__30957\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__30974\,
            I => \N__30957\
        );

    \I__5793\ : Sp12to4
    port map (
            O => \N__30971\,
            I => \N__30954\
        );

    \I__5792\ : LocalMux
    port map (
            O => \N__30968\,
            I => \N__30951\
        );

    \I__5791\ : Span12Mux_v
    port map (
            O => \N__30965\,
            I => \N__30948\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__30962\,
            I => \N__30945\
        );

    \I__5789\ : Span4Mux_v
    port map (
            O => \N__30957\,
            I => \N__30942\
        );

    \I__5788\ : Span12Mux_h
    port map (
            O => \N__30954\,
            I => \N__30939\
        );

    \I__5787\ : Span12Mux_s6_h
    port map (
            O => \N__30951\,
            I => \N__30936\
        );

    \I__5786\ : Span12Mux_v
    port map (
            O => \N__30948\,
            I => \N__30933\
        );

    \I__5785\ : Span12Mux_h
    port map (
            O => \N__30945\,
            I => \N__30930\
        );

    \I__5784\ : Span4Mux_h
    port map (
            O => \N__30942\,
            I => \N__30927\
        );

    \I__5783\ : Span12Mux_v
    port map (
            O => \N__30939\,
            I => \N__30922\
        );

    \I__5782\ : Span12Mux_h
    port map (
            O => \N__30936\,
            I => \N__30922\
        );

    \I__5781\ : Span12Mux_h
    port map (
            O => \N__30933\,
            I => \N__30917\
        );

    \I__5780\ : Span12Mux_v
    port map (
            O => \N__30930\,
            I => \N__30917\
        );

    \I__5779\ : Span4Mux_v
    port map (
            O => \N__30927\,
            I => \N__30914\
        );

    \I__5778\ : Odrv12
    port map (
            O => \N__30922\,
            I => start_stop_c
        );

    \I__5777\ : Odrv12
    port map (
            O => \N__30917\,
            I => start_stop_c
        );

    \I__5776\ : Odrv4
    port map (
            O => \N__30914\,
            I => start_stop_c
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__30907\,
            I => \N__30902\
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__30906\,
            I => \N__30899\
        );

    \I__5773\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30896\
        );

    \I__5772\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30891\
        );

    \I__5771\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30891\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__30896\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__30891\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__5768\ : InMux
    port map (
            O => \N__30886\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__5767\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30878\
        );

    \I__5766\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30875\
        );

    \I__5765\ : InMux
    port map (
            O => \N__30881\,
            I => \N__30872\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__30878\,
            I => \N__30869\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__30875\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__30872\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__30869\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__5760\ : InMux
    port map (
            O => \N__30862\,
            I => \bfn_13_9_0_\
        );

    \I__5759\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30854\
        );

    \I__5758\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30851\
        );

    \I__5757\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30848\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__30854\,
            I => \N__30845\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__30851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__30848\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__5753\ : Odrv4
    port map (
            O => \N__30845\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__5752\ : InMux
    port map (
            O => \N__30838\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__30835\,
            I => \N__30830\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__30834\,
            I => \N__30827\
        );

    \I__5749\ : InMux
    port map (
            O => \N__30833\,
            I => \N__30824\
        );

    \I__5748\ : InMux
    port map (
            O => \N__30830\,
            I => \N__30819\
        );

    \I__5747\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30819\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__30824\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__30819\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__5744\ : InMux
    port map (
            O => \N__30814\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__30811\,
            I => \N__30806\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__30810\,
            I => \N__30803\
        );

    \I__5741\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30800\
        );

    \I__5740\ : InMux
    port map (
            O => \N__30806\,
            I => \N__30795\
        );

    \I__5739\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30795\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__30800\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__30795\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30790\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__5735\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30782\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30777\
        );

    \I__5733\ : InMux
    port map (
            O => \N__30785\,
            I => \N__30777\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__30782\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__30777\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__5730\ : InMux
    port map (
            O => \N__30772\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__5729\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30764\
        );

    \I__5728\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30759\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30767\,
            I => \N__30759\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__30764\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__30759\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__5724\ : InMux
    port map (
            O => \N__30754\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__30751\,
            I => \N__30746\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__30750\,
            I => \N__30743\
        );

    \I__5721\ : InMux
    port map (
            O => \N__30749\,
            I => \N__30740\
        );

    \I__5720\ : InMux
    port map (
            O => \N__30746\,
            I => \N__30735\
        );

    \I__5719\ : InMux
    port map (
            O => \N__30743\,
            I => \N__30735\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__30740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__30735\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30730\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__30727\,
            I => \N__30722\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__30726\,
            I => \N__30719\
        );

    \I__5713\ : InMux
    port map (
            O => \N__30725\,
            I => \N__30716\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30711\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30711\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__30716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__30711\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__5708\ : InMux
    port map (
            O => \N__30706\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__5707\ : CascadeMux
    port map (
            O => \N__30703\,
            I => \N__30698\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__30702\,
            I => \N__30695\
        );

    \I__5705\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30692\
        );

    \I__5704\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30687\
        );

    \I__5703\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30687\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__30692\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__30687\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__5700\ : InMux
    port map (
            O => \N__30682\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__5699\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30674\
        );

    \I__5698\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30671\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30677\,
            I => \N__30668\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__30674\,
            I => \N__30665\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__30671\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30668\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5693\ : Odrv4
    port map (
            O => \N__30665\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30658\,
            I => \bfn_13_8_0_\
        );

    \I__5691\ : InMux
    port map (
            O => \N__30655\,
            I => \N__30650\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30647\
        );

    \I__5689\ : InMux
    port map (
            O => \N__30653\,
            I => \N__30644\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__30650\,
            I => \N__30641\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__30647\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__30644\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__30641\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__5684\ : InMux
    port map (
            O => \N__30634\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__30631\,
            I => \N__30626\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__30630\,
            I => \N__30623\
        );

    \I__5681\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30620\
        );

    \I__5680\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30615\
        );

    \I__5679\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30615\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__30620\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__30615\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__5676\ : InMux
    port map (
            O => \N__30610\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__5675\ : CascadeMux
    port map (
            O => \N__30607\,
            I => \N__30602\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__30606\,
            I => \N__30599\
        );

    \I__5673\ : InMux
    port map (
            O => \N__30605\,
            I => \N__30596\
        );

    \I__5672\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30591\
        );

    \I__5671\ : InMux
    port map (
            O => \N__30599\,
            I => \N__30591\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__30596\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__30591\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30586\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__5667\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30578\
        );

    \I__5666\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30573\
        );

    \I__5665\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30573\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__30578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__30573\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__5662\ : InMux
    port map (
            O => \N__30568\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30560\
        );

    \I__5660\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30555\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30555\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__30560\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__30555\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30550\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__5655\ : CascadeMux
    port map (
            O => \N__30547\,
            I => \N__30542\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__30546\,
            I => \N__30539\
        );

    \I__5653\ : InMux
    port map (
            O => \N__30545\,
            I => \N__30536\
        );

    \I__5652\ : InMux
    port map (
            O => \N__30542\,
            I => \N__30531\
        );

    \I__5651\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30531\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__30536\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__30531\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__5648\ : InMux
    port map (
            O => \N__30526\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__5647\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30520\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30520\,
            I => \N__30516\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__30519\,
            I => \N__30512\
        );

    \I__5644\ : Span4Mux_v
    port map (
            O => \N__30516\,
            I => \N__30508\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30505\
        );

    \I__5642\ : InMux
    port map (
            O => \N__30512\,
            I => \N__30502\
        );

    \I__5641\ : InMux
    port map (
            O => \N__30511\,
            I => \N__30499\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__30508\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__30505\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__30502\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30499\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__5636\ : InMux
    port map (
            O => \N__30490\,
            I => \N__30487\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__30487\,
            I => \N__30477\
        );

    \I__5634\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30474\
        );

    \I__5633\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30469\
        );

    \I__5632\ : InMux
    port map (
            O => \N__30484\,
            I => \N__30469\
        );

    \I__5631\ : InMux
    port map (
            O => \N__30483\,
            I => \N__30460\
        );

    \I__5630\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30460\
        );

    \I__5629\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30460\
        );

    \I__5628\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30457\
        );

    \I__5627\ : Span4Mux_v
    port map (
            O => \N__30477\,
            I => \N__30452\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__30474\,
            I => \N__30449\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__30469\,
            I => \N__30446\
        );

    \I__5624\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30441\
        );

    \I__5623\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30441\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__30460\,
            I => \N__30438\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__30457\,
            I => \N__30434\
        );

    \I__5620\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30429\
        );

    \I__5619\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30429\
        );

    \I__5618\ : Span4Mux_v
    port map (
            O => \N__30452\,
            I => \N__30411\
        );

    \I__5617\ : Span4Mux_v
    port map (
            O => \N__30449\,
            I => \N__30411\
        );

    \I__5616\ : Span4Mux_v
    port map (
            O => \N__30446\,
            I => \N__30411\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30408\
        );

    \I__5614\ : Span4Mux_h
    port map (
            O => \N__30438\,
            I => \N__30405\
        );

    \I__5613\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30402\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__30434\,
            I => \N__30397\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30429\,
            I => \N__30397\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30382\
        );

    \I__5609\ : InMux
    port map (
            O => \N__30427\,
            I => \N__30382\
        );

    \I__5608\ : InMux
    port map (
            O => \N__30426\,
            I => \N__30382\
        );

    \I__5607\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30382\
        );

    \I__5606\ : InMux
    port map (
            O => \N__30424\,
            I => \N__30382\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30382\
        );

    \I__5604\ : InMux
    port map (
            O => \N__30422\,
            I => \N__30382\
        );

    \I__5603\ : InMux
    port map (
            O => \N__30421\,
            I => \N__30373\
        );

    \I__5602\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30373\
        );

    \I__5601\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30373\
        );

    \I__5600\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30373\
        );

    \I__5599\ : Odrv4
    port map (
            O => \N__30411\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__30408\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5597\ : Odrv4
    port map (
            O => \N__30405\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__30402\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__30397\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__30382\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__30373\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__5592\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30353\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30357\,
            I => \N__30350\
        );

    \I__5590\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30347\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30344\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__30350\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__30347\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__5586\ : Odrv12
    port map (
            O => \N__30344\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30337\,
            I => \N__30332\
        );

    \I__5584\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30329\
        );

    \I__5583\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30326\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__30332\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__30329\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__30326\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__5579\ : InMux
    port map (
            O => \N__30319\,
            I => \bfn_13_7_0_\
        );

    \I__5578\ : InMux
    port map (
            O => \N__30316\,
            I => \N__30311\
        );

    \I__5577\ : InMux
    port map (
            O => \N__30315\,
            I => \N__30308\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30314\,
            I => \N__30305\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__30311\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__30308\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__30305\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__5572\ : InMux
    port map (
            O => \N__30298\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__5571\ : CascadeMux
    port map (
            O => \N__30295\,
            I => \N__30290\
        );

    \I__5570\ : CascadeMux
    port map (
            O => \N__30294\,
            I => \N__30287\
        );

    \I__5569\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30284\
        );

    \I__5568\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30279\
        );

    \I__5567\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30279\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__30284\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__30279\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__5564\ : InMux
    port map (
            O => \N__30274\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__30271\,
            I => \N__30266\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__30270\,
            I => \N__30263\
        );

    \I__5561\ : InMux
    port map (
            O => \N__30269\,
            I => \N__30260\
        );

    \I__5560\ : InMux
    port map (
            O => \N__30266\,
            I => \N__30255\
        );

    \I__5559\ : InMux
    port map (
            O => \N__30263\,
            I => \N__30255\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__30260\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__30255\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__5556\ : InMux
    port map (
            O => \N__30250\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30247\,
            I => \N__30242\
        );

    \I__5554\ : InMux
    port map (
            O => \N__30246\,
            I => \N__30237\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30245\,
            I => \N__30237\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__30242\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__30237\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30232\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__5549\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30224\
        );

    \I__5548\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30219\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30219\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30224\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__30219\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__5544\ : InMux
    port map (
            O => \N__30214\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__5543\ : InMux
    port map (
            O => \N__30211\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30208\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30205\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__5540\ : InMux
    port map (
            O => \N__30202\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__30199\,
            I => \N__30196\
        );

    \I__5538\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30193\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__30193\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__5536\ : InMux
    port map (
            O => \N__30190\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__5535\ : InMux
    port map (
            O => \N__30187\,
            I => \bfn_12_26_0_\
        );

    \I__5534\ : InMux
    port map (
            O => \N__30184\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__5533\ : InMux
    port map (
            O => \N__30181\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30178\,
            I => \N__30175\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__30175\,
            I => \N__30169\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30166\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30163\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30172\,
            I => \N__30160\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__30169\,
            I => \N__30157\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__30166\,
            I => \N__30154\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__30163\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30160\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__30157\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5522\ : Odrv4
    port map (
            O => \N__30154\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30142\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__30142\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__5519\ : InMux
    port map (
            O => \N__30139\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30136\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30133\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__5516\ : InMux
    port map (
            O => \N__30130\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__5515\ : InMux
    port map (
            O => \N__30127\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30121\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30118\
        );

    \I__5512\ : Odrv12
    port map (
            O => \N__30118\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30115\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__5510\ : InMux
    port map (
            O => \N__30112\,
            I => \N__30109\
        );

    \I__5509\ : LocalMux
    port map (
            O => \N__30109\,
            I => \N__30106\
        );

    \I__5508\ : Odrv12
    port map (
            O => \N__30106\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30103\,
            I => \bfn_12_25_0_\
        );

    \I__5506\ : InMux
    port map (
            O => \N__30100\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__5505\ : InMux
    port map (
            O => \N__30097\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__5504\ : CascadeMux
    port map (
            O => \N__30094\,
            I => \N__30090\
        );

    \I__5503\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30087\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30084\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__30087\,
            I => \current_shift_inst.z_i_31\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__30084\,
            I => \current_shift_inst.z_i_31\
        );

    \I__5499\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30076\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__30076\,
            I => \N__30073\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__30073\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\
        );

    \I__5496\ : IoInMux
    port map (
            O => \N__30070\,
            I => \N__30067\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__30067\,
            I => \N__30064\
        );

    \I__5494\ : Span4Mux_s2_v
    port map (
            O => \N__30064\,
            I => \N__30061\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__30061\,
            I => \N__30058\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__30058\,
            I => \current_shift_inst.timer_phase.N_188_i\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30052\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30052\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__5489\ : InMux
    port map (
            O => \N__30049\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__5488\ : IoInMux
    port map (
            O => \N__30046\,
            I => \N__30043\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30043\,
            I => \N__30040\
        );

    \I__5486\ : Span4Mux_s3_v
    port map (
            O => \N__30040\,
            I => \N__30037\
        );

    \I__5485\ : Span4Mux_h
    port map (
            O => \N__30037\,
            I => \N__30034\
        );

    \I__5484\ : Sp12to4
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__5483\ : Span12Mux_v
    port map (
            O => \N__30031\,
            I => \N__30027\
        );

    \I__5482\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30024\
        );

    \I__5481\ : Odrv12
    port map (
            O => \N__30027\,
            I => s1_phy_c
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30024\,
            I => s1_phy_c
        );

    \I__5479\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30016\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30016\,
            I => \N__30013\
        );

    \I__5477\ : Span4Mux_v
    port map (
            O => \N__30013\,
            I => \N__30010\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__30010\,
            I => \N__30007\
        );

    \I__5475\ : Odrv4
    port map (
            O => \N__30007\,
            I => \phase_controller_inst1.stoper_tr.N_21\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30004\,
            I => \N__30001\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__30001\,
            I => \N__29998\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__29998\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3\
        );

    \I__5471\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29992\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__29992\,
            I => \N__29987\
        );

    \I__5469\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29982\
        );

    \I__5468\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29982\
        );

    \I__5467\ : Odrv4
    port map (
            O => \N__29987\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__29982\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__5465\ : InMux
    port map (
            O => \N__29977\,
            I => \N__29974\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__29974\,
            I => \N__29971\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__29971\,
            I => \N__29965\
        );

    \I__5462\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29962\
        );

    \I__5461\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29959\
        );

    \I__5460\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29956\
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__29965\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__29962\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__29959\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__29956\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__29947\,
            I => \N__29943\
        );

    \I__5454\ : InMux
    port map (
            O => \N__29946\,
            I => \N__29940\
        );

    \I__5453\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29937\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29933\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__29937\,
            I => \N__29930\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__29936\,
            I => \N__29927\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__29933\,
            I => \N__29923\
        );

    \I__5448\ : Span4Mux_h
    port map (
            O => \N__29930\,
            I => \N__29920\
        );

    \I__5447\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29917\
        );

    \I__5446\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29914\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__29923\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5444\ : Odrv4
    port map (
            O => \N__29920\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__29917\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__29914\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__5441\ : InMux
    port map (
            O => \N__29905\,
            I => \N__29900\
        );

    \I__5440\ : InMux
    port map (
            O => \N__29904\,
            I => \N__29897\
        );

    \I__5439\ : InMux
    port map (
            O => \N__29903\,
            I => \N__29894\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__29900\,
            I => \N__29891\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__29897\,
            I => \N__29886\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__29894\,
            I => \N__29886\
        );

    \I__5435\ : Odrv4
    port map (
            O => \N__29891\,
            I => \il_min_comp1_D2\
        );

    \I__5434\ : Odrv4
    port map (
            O => \N__29886\,
            I => \il_min_comp1_D2\
        );

    \I__5433\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29874\
        );

    \I__5432\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29871\
        );

    \I__5431\ : CascadeMux
    port map (
            O => \N__29879\,
            I => \N__29868\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__29878\,
            I => \N__29865\
        );

    \I__5429\ : CascadeMux
    port map (
            O => \N__29877\,
            I => \N__29862\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29857\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__29871\,
            I => \N__29857\
        );

    \I__5426\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29854\
        );

    \I__5425\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29851\
        );

    \I__5424\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29848\
        );

    \I__5423\ : Span12Mux_v
    port map (
            O => \N__29857\,
            I => \N__29845\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__29854\,
            I => \N__29840\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__29851\,
            I => \N__29840\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__29848\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5419\ : Odrv12
    port map (
            O => \N__29845\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5418\ : Odrv4
    port map (
            O => \N__29840\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__5417\ : InMux
    port map (
            O => \N__29833\,
            I => \N__29829\
        );

    \I__5416\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29826\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__29829\,
            I => \N__29823\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__29826\,
            I => \N__29819\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__29823\,
            I => \N__29816\
        );

    \I__5412\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29812\
        );

    \I__5411\ : Span4Mux_h
    port map (
            O => \N__29819\,
            I => \N__29807\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__29816\,
            I => \N__29807\
        );

    \I__5409\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29804\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__29812\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__29807\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__29804\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__5405\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29794\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__29794\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__5403\ : InMux
    port map (
            O => \N__29791\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__5402\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29785\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__29785\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__5400\ : InMux
    port map (
            O => \N__29782\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__29779\,
            I => \N__29776\
        );

    \I__5398\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29773\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__29773\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29770\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__5395\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29764\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__29764\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__5393\ : InMux
    port map (
            O => \N__29761\,
            I => \bfn_12_10_0_\
        );

    \I__5392\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29755\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__29755\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__5390\ : InMux
    port map (
            O => \N__29752\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__5389\ : InMux
    port map (
            O => \N__29749\,
            I => \N__29746\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__29746\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__5387\ : InMux
    port map (
            O => \N__29743\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__29740\,
            I => \N__29737\
        );

    \I__5385\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29734\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__29734\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29731\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29728\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__29725\,
            I => \N__29722\
        );

    \I__5380\ : InMux
    port map (
            O => \N__29722\,
            I => \N__29715\
        );

    \I__5379\ : InMux
    port map (
            O => \N__29721\,
            I => \N__29715\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__29720\,
            I => \N__29712\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29709\
        );

    \I__5376\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29706\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__29709\,
            I => \N__29703\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__29706\,
            I => \N__29700\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__29703\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__29700\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__5371\ : CEMux
    port map (
            O => \N__29695\,
            I => \N__29680\
        );

    \I__5370\ : CEMux
    port map (
            O => \N__29694\,
            I => \N__29680\
        );

    \I__5369\ : CEMux
    port map (
            O => \N__29693\,
            I => \N__29680\
        );

    \I__5368\ : CEMux
    port map (
            O => \N__29692\,
            I => \N__29680\
        );

    \I__5367\ : CEMux
    port map (
            O => \N__29691\,
            I => \N__29680\
        );

    \I__5366\ : GlobalMux
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__5365\ : gio2CtrlBuf
    port map (
            O => \N__29677\,
            I => \delay_measurement_inst.delay_hc_timer.N_336_i_g\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29674\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__5363\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29668\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29665\
        );

    \I__5361\ : Span4Mux_h
    port map (
            O => \N__29665\,
            I => \N__29660\
        );

    \I__5360\ : InMux
    port map (
            O => \N__29664\,
            I => \N__29657\
        );

    \I__5359\ : InMux
    port map (
            O => \N__29663\,
            I => \N__29654\
        );

    \I__5358\ : Odrv4
    port map (
            O => \N__29660\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__29657\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__29654\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29647\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29641\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29638\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__29638\,
            I => \N__29633\
        );

    \I__5351\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29630\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29627\
        );

    \I__5349\ : Odrv4
    port map (
            O => \N__29633\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29630\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__29627\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__5346\ : InMux
    port map (
            O => \N__29620\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__5345\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29612\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29609\
        );

    \I__5343\ : CascadeMux
    port map (
            O => \N__29615\,
            I => \N__29606\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__29612\,
            I => \N__29603\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29600\
        );

    \I__5340\ : InMux
    port map (
            O => \N__29606\,
            I => \N__29597\
        );

    \I__5339\ : Odrv12
    port map (
            O => \N__29603\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__29600\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__29597\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__5336\ : InMux
    port map (
            O => \N__29590\,
            I => \bfn_12_9_0_\
        );

    \I__5335\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29583\
        );

    \I__5334\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29580\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__29583\,
            I => \N__29577\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__29580\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5331\ : Odrv4
    port map (
            O => \N__29577\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__5330\ : InMux
    port map (
            O => \N__29572\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__5329\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29563\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29563\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29563\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__5326\ : InMux
    port map (
            O => \N__29560\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__29557\,
            I => \N__29554\
        );

    \I__5324\ : InMux
    port map (
            O => \N__29554\,
            I => \N__29548\
        );

    \I__5323\ : InMux
    port map (
            O => \N__29553\,
            I => \N__29548\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__29548\,
            I => \N__29545\
        );

    \I__5321\ : Odrv4
    port map (
            O => \N__29545\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__5320\ : InMux
    port map (
            O => \N__29542\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__5319\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29536\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__29536\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__5317\ : InMux
    port map (
            O => \N__29533\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__5316\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29525\
        );

    \I__5315\ : InMux
    port map (
            O => \N__29529\,
            I => \N__29522\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29528\,
            I => \N__29519\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29525\,
            I => \N__29512\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__29522\,
            I => \N__29512\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__29519\,
            I => \N__29512\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__29512\,
            I => \N__29508\
        );

    \I__5309\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29505\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__29508\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__29505\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__5306\ : InMux
    port map (
            O => \N__29500\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__29497\,
            I => \N__29492\
        );

    \I__5304\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29489\
        );

    \I__5303\ : InMux
    port map (
            O => \N__29495\,
            I => \N__29486\
        );

    \I__5302\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29483\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__29489\,
            I => \N__29476\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__29486\,
            I => \N__29476\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__29483\,
            I => \N__29476\
        );

    \I__5298\ : Span4Mux_v
    port map (
            O => \N__29476\,
            I => \N__29472\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29469\
        );

    \I__5296\ : Odrv4
    port map (
            O => \N__29472\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__29469\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29464\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__5293\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29458\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__29458\,
            I => \N__29453\
        );

    \I__5291\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29450\
        );

    \I__5290\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29447\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__29453\,
            I => \N__29442\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29442\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__29447\,
            I => \N__29439\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__29442\,
            I => \N__29435\
        );

    \I__5285\ : Span4Mux_h
    port map (
            O => \N__29439\,
            I => \N__29432\
        );

    \I__5284\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29429\
        );

    \I__5283\ : Odrv4
    port map (
            O => \N__29435\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__29432\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__29429\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__5280\ : InMux
    port map (
            O => \N__29422\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__29419\,
            I => \N__29416\
        );

    \I__5278\ : InMux
    port map (
            O => \N__29416\,
            I => \N__29412\
        );

    \I__5277\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29409\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29406\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__29409\,
            I => \N__29402\
        );

    \I__5274\ : Span4Mux_h
    port map (
            O => \N__29406\,
            I => \N__29399\
        );

    \I__5273\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29396\
        );

    \I__5272\ : Span4Mux_h
    port map (
            O => \N__29402\,
            I => \N__29393\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__29399\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__29396\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__29393\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__5268\ : InMux
    port map (
            O => \N__29386\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__5267\ : InMux
    port map (
            O => \N__29383\,
            I => \N__29380\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__29380\,
            I => \N__29376\
        );

    \I__5265\ : InMux
    port map (
            O => \N__29379\,
            I => \N__29373\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__29376\,
            I => \N__29369\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__29373\,
            I => \N__29366\
        );

    \I__5262\ : InMux
    port map (
            O => \N__29372\,
            I => \N__29363\
        );

    \I__5261\ : Odrv4
    port map (
            O => \N__29369\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__29366\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__29363\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__5258\ : InMux
    port map (
            O => \N__29356\,
            I => \bfn_12_8_0_\
        );

    \I__5257\ : CascadeMux
    port map (
            O => \N__29353\,
            I => \N__29349\
        );

    \I__5256\ : CascadeMux
    port map (
            O => \N__29352\,
            I => \N__29345\
        );

    \I__5255\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29342\
        );

    \I__5254\ : InMux
    port map (
            O => \N__29348\,
            I => \N__29339\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29336\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__29342\,
            I => \N__29333\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__29339\,
            I => \N__29330\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__29336\,
            I => \N__29327\
        );

    \I__5249\ : Span4Mux_h
    port map (
            O => \N__29333\,
            I => \N__29324\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__29330\,
            I => \N__29319\
        );

    \I__5247\ : Span4Mux_h
    port map (
            O => \N__29327\,
            I => \N__29319\
        );

    \I__5246\ : Odrv4
    port map (
            O => \N__29324\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__29319\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__5244\ : InMux
    port map (
            O => \N__29314\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__5243\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29308\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29303\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29300\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__29306\,
            I => \N__29297\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__29303\,
            I => \N__29294\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__29300\,
            I => \N__29291\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29288\
        );

    \I__5236\ : Odrv4
    port map (
            O => \N__29294\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__29291\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__29288\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29281\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__5232\ : InMux
    port map (
            O => \N__29278\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__5231\ : InMux
    port map (
            O => \N__29275\,
            I => \N__29272\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__29272\,
            I => \N__29263\
        );

    \I__5229\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29260\
        );

    \I__5228\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29255\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29255\
        );

    \I__5226\ : InMux
    port map (
            O => \N__29268\,
            I => \N__29252\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29247\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29266\,
            I => \N__29247\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__29263\,
            I => \N__29240\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29260\,
            I => \N__29240\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__29255\,
            I => \N__29240\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__29252\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__29247\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__29240\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29233\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__29230\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29227\,
            I => \N__29223\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29220\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__29223\,
            I => \N__29215\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__29220\,
            I => \N__29215\
        );

    \I__5211\ : Span4Mux_v
    port map (
            O => \N__29215\,
            I => \N__29212\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__29212\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__5209\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29205\
        );

    \I__5208\ : CascadeMux
    port map (
            O => \N__29208\,
            I => \N__29201\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29205\,
            I => \N__29198\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29195\
        );

    \I__5205\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29192\
        );

    \I__5204\ : Span4Mux_v
    port map (
            O => \N__29198\,
            I => \N__29187\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29187\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__29192\,
            I => \N__29182\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__29187\,
            I => \N__29182\
        );

    \I__5200\ : Odrv4
    port map (
            O => \N__29182\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29179\,
            I => \N__29175\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29172\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29175\,
            I => \N__29168\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__29172\,
            I => \N__29165\
        );

    \I__5195\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29162\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__29168\,
            I => \N__29159\
        );

    \I__5193\ : Odrv12
    port map (
            O => \N__29165\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__29162\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__5191\ : Odrv4
    port map (
            O => \N__29159\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29152\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__5189\ : CascadeMux
    port map (
            O => \N__29149\,
            I => \N__29145\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29141\
        );

    \I__5187\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29138\
        );

    \I__5186\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29135\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29130\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__29138\,
            I => \N__29130\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29135\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__29130\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29125\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__5180\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29118\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__29121\,
            I => \N__29114\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29111\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29106\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29114\,
            I => \N__29106\
        );

    \I__5175\ : Span4Mux_h
    port map (
            O => \N__29111\,
            I => \N__29101\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__29106\,
            I => \N__29101\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__29101\,
            I => \N__29097\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29094\
        );

    \I__5171\ : Odrv4
    port map (
            O => \N__29097\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__29094\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__5169\ : InMux
    port map (
            O => \N__29089\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__5168\ : CascadeMux
    port map (
            O => \N__29086\,
            I => \N__29083\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29083\,
            I => \N__29080\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29077\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__29077\,
            I => \current_shift_inst.control_input_1_axb_22\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29070\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__29073\,
            I => \N__29067\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__29070\,
            I => \N__29064\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29061\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__29064\,
            I => \N__29056\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__29061\,
            I => \N__29056\
        );

    \I__5158\ : Span4Mux_h
    port map (
            O => \N__29056\,
            I => \N__29053\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__29053\,
            I => \N__29050\
        );

    \I__5156\ : Odrv4
    port map (
            O => \N__29050\,
            I => \current_shift_inst.control_inputZ0Z_22\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29047\,
            I => \current_shift_inst.control_input_1_cry_21\
        );

    \I__5154\ : CascadeMux
    port map (
            O => \N__29044\,
            I => \N__29041\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29041\,
            I => \N__29038\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__29038\,
            I => \N__29035\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__29035\,
            I => \current_shift_inst.control_input_1_axb_23\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29028\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__29031\,
            I => \N__29025\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__29028\,
            I => \N__29022\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29025\,
            I => \N__29019\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__29022\,
            I => \N__29016\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__29019\,
            I => \N__29013\
        );

    \I__5144\ : Span4Mux_h
    port map (
            O => \N__29016\,
            I => \N__29008\
        );

    \I__5143\ : Span4Mux_v
    port map (
            O => \N__29013\,
            I => \N__29008\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__29008\,
            I => \current_shift_inst.control_inputZ0Z_23\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29005\,
            I => \current_shift_inst.control_input_1_cry_22\
        );

    \I__5140\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28999\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__28999\,
            I => \current_shift_inst.control_input_1_axb_24\
        );

    \I__5138\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28992\
        );

    \I__5137\ : CascadeMux
    port map (
            O => \N__28995\,
            I => \N__28989\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__28992\,
            I => \N__28986\
        );

    \I__5135\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28983\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__28986\,
            I => \N__28978\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__28983\,
            I => \N__28978\
        );

    \I__5132\ : Span4Mux_h
    port map (
            O => \N__28978\,
            I => \N__28975\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__28975\,
            I => \current_shift_inst.control_inputZ0Z_24\
        );

    \I__5130\ : InMux
    port map (
            O => \N__28972\,
            I => \bfn_11_23_0_\
        );

    \I__5129\ : CEMux
    port map (
            O => \N__28969\,
            I => \N__28966\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28960\
        );

    \I__5127\ : CEMux
    port map (
            O => \N__28965\,
            I => \N__28957\
        );

    \I__5126\ : CEMux
    port map (
            O => \N__28964\,
            I => \N__28954\
        );

    \I__5125\ : CEMux
    port map (
            O => \N__28963\,
            I => \N__28951\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__28960\,
            I => \N__28945\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28945\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28942\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28939\
        );

    \I__5120\ : CEMux
    port map (
            O => \N__28950\,
            I => \N__28936\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__28945\,
            I => \N__28933\
        );

    \I__5118\ : Span4Mux_v
    port map (
            O => \N__28942\,
            I => \N__28930\
        );

    \I__5117\ : Span4Mux_v
    port map (
            O => \N__28939\,
            I => \N__28927\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28924\
        );

    \I__5115\ : Span4Mux_h
    port map (
            O => \N__28933\,
            I => \N__28921\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__28930\,
            I => \N__28918\
        );

    \I__5113\ : Sp12to4
    port map (
            O => \N__28927\,
            I => \N__28915\
        );

    \I__5112\ : Span4Mux_v
    port map (
            O => \N__28924\,
            I => \N__28912\
        );

    \I__5111\ : Span4Mux_h
    port map (
            O => \N__28921\,
            I => \N__28909\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__28918\,
            I => \N__28906\
        );

    \I__5109\ : Span12Mux_h
    port map (
            O => \N__28915\,
            I => \N__28903\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__28912\,
            I => \N__28900\
        );

    \I__5107\ : Span4Mux_v
    port map (
            O => \N__28909\,
            I => \N__28897\
        );

    \I__5106\ : Span4Mux_v
    port map (
            O => \N__28906\,
            I => \N__28894\
        );

    \I__5105\ : Span12Mux_v
    port map (
            O => \N__28903\,
            I => \N__28889\
        );

    \I__5104\ : Sp12to4
    port map (
            O => \N__28900\,
            I => \N__28889\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__28897\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__28894\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__5101\ : Odrv12
    port map (
            O => \N__28889\,
            I => \current_shift_inst.phase_valid_RNISLORZ0Z2\
        );

    \I__5100\ : InMux
    port map (
            O => \N__28882\,
            I => \current_shift_inst.control_input_1_cry_24\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__28879\,
            I => \N__28876\
        );

    \I__5098\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28873\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28870\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__28870\,
            I => \current_shift_inst.control_input_1_cry_24_THRU_CO\
        );

    \I__5095\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28863\
        );

    \I__5094\ : CascadeMux
    port map (
            O => \N__28866\,
            I => \N__28860\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__28863\,
            I => \N__28857\
        );

    \I__5092\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28854\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__28857\,
            I => \N__28849\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__28854\,
            I => \N__28849\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__28849\,
            I => \N__28846\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__28846\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\
        );

    \I__5087\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28840\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__28840\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\
        );

    \I__5085\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28834\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__28834\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\
        );

    \I__5083\ : CascadeMux
    port map (
            O => \N__28831\,
            I => \N__28828\
        );

    \I__5082\ : InMux
    port map (
            O => \N__28828\,
            I => \N__28825\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__28825\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__28822\,
            I => \N__28819\
        );

    \I__5079\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28816\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__28816\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__28813\,
            I => \N__28810\
        );

    \I__5076\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28807\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__28807\,
            I => \N__28804\
        );

    \I__5074\ : Odrv4
    port map (
            O => \N__28804\,
            I => \current_shift_inst.control_input_1_axb_14\
        );

    \I__5073\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28797\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__28800\,
            I => \N__28794\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28791\
        );

    \I__5070\ : InMux
    port map (
            O => \N__28794\,
            I => \N__28788\
        );

    \I__5069\ : Span4Mux_h
    port map (
            O => \N__28791\,
            I => \N__28783\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28783\
        );

    \I__5067\ : Span4Mux_h
    port map (
            O => \N__28783\,
            I => \N__28780\
        );

    \I__5066\ : Odrv4
    port map (
            O => \N__28780\,
            I => \current_shift_inst.control_inputZ0Z_14\
        );

    \I__5065\ : InMux
    port map (
            O => \N__28777\,
            I => \current_shift_inst.control_input_1_cry_13\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__28774\,
            I => \N__28771\
        );

    \I__5063\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28768\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__28768\,
            I => \N__28765\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__28765\,
            I => \current_shift_inst.control_input_1_axb_15\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28758\
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__28761\,
            I => \N__28755\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__28758\,
            I => \N__28752\
        );

    \I__5057\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28749\
        );

    \I__5056\ : Span4Mux_v
    port map (
            O => \N__28752\,
            I => \N__28746\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__28749\,
            I => \N__28743\
        );

    \I__5054\ : Sp12to4
    port map (
            O => \N__28746\,
            I => \N__28740\
        );

    \I__5053\ : Span4Mux_v
    port map (
            O => \N__28743\,
            I => \N__28737\
        );

    \I__5052\ : Odrv12
    port map (
            O => \N__28740\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__28737\,
            I => \current_shift_inst.control_inputZ0Z_15\
        );

    \I__5050\ : InMux
    port map (
            O => \N__28732\,
            I => \current_shift_inst.control_input_1_cry_14\
        );

    \I__5049\ : InMux
    port map (
            O => \N__28729\,
            I => \N__28726\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__28726\,
            I => \current_shift_inst.control_input_1_axb_16\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28723\,
            I => \N__28719\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__28722\,
            I => \N__28716\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__28719\,
            I => \N__28713\
        );

    \I__5044\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28710\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__28713\,
            I => \N__28707\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__28710\,
            I => \N__28704\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__28707\,
            I => \N__28699\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__28704\,
            I => \N__28699\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__28699\,
            I => \current_shift_inst.control_inputZ0Z_16\
        );

    \I__5038\ : InMux
    port map (
            O => \N__28696\,
            I => \bfn_11_22_0_\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__28690\,
            I => \N__28687\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__28687\,
            I => \current_shift_inst.control_input_1_axb_17\
        );

    \I__5034\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28680\
        );

    \I__5033\ : InMux
    port map (
            O => \N__28683\,
            I => \N__28677\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28674\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__28677\,
            I => \N__28671\
        );

    \I__5030\ : Span12Mux_s11_h
    port map (
            O => \N__28674\,
            I => \N__28668\
        );

    \I__5029\ : Span4Mux_h
    port map (
            O => \N__28671\,
            I => \N__28665\
        );

    \I__5028\ : Odrv12
    port map (
            O => \N__28668\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__28665\,
            I => \current_shift_inst.control_inputZ0Z_17\
        );

    \I__5026\ : InMux
    port map (
            O => \N__28660\,
            I => \current_shift_inst.control_input_1_cry_16\
        );

    \I__5025\ : InMux
    port map (
            O => \N__28657\,
            I => \N__28654\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__28654\,
            I => \N__28651\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__28651\,
            I => \current_shift_inst.control_input_1_axb_18\
        );

    \I__5022\ : CascadeMux
    port map (
            O => \N__28648\,
            I => \N__28644\
        );

    \I__5021\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28641\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28638\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__28641\,
            I => \N__28635\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__28638\,
            I => \N__28632\
        );

    \I__5017\ : Span4Mux_h
    port map (
            O => \N__28635\,
            I => \N__28627\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__28632\,
            I => \N__28627\
        );

    \I__5015\ : Odrv4
    port map (
            O => \N__28627\,
            I => \current_shift_inst.control_inputZ0Z_18\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28624\,
            I => \current_shift_inst.control_input_1_cry_17\
        );

    \I__5013\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28615\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__28615\,
            I => \current_shift_inst.control_input_1_axb_19\
        );

    \I__5010\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28608\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__28611\,
            I => \N__28605\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28602\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28599\
        );

    \I__5006\ : Span4Mux_h
    port map (
            O => \N__28602\,
            I => \N__28594\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28594\
        );

    \I__5004\ : Span4Mux_h
    port map (
            O => \N__28594\,
            I => \N__28591\
        );

    \I__5003\ : Odrv4
    port map (
            O => \N__28591\,
            I => \current_shift_inst.control_inputZ0Z_19\
        );

    \I__5002\ : InMux
    port map (
            O => \N__28588\,
            I => \current_shift_inst.control_input_1_cry_18\
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__5000\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28579\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__28579\,
            I => \N__28576\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__28576\,
            I => \current_shift_inst.control_input_1_axb_20\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__28573\,
            I => \N__28569\
        );

    \I__4996\ : InMux
    port map (
            O => \N__28572\,
            I => \N__28566\
        );

    \I__4995\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28563\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28558\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28558\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__28558\,
            I => \N__28555\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__28555\,
            I => \current_shift_inst.control_inputZ0Z_20\
        );

    \I__4990\ : InMux
    port map (
            O => \N__28552\,
            I => \current_shift_inst.control_input_1_cry_19\
        );

    \I__4989\ : CascadeMux
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__4988\ : InMux
    port map (
            O => \N__28546\,
            I => \N__28543\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__28543\,
            I => \N__28540\
        );

    \I__4986\ : Odrv4
    port map (
            O => \N__28540\,
            I => \current_shift_inst.control_input_1_axb_21\
        );

    \I__4985\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28533\
        );

    \I__4984\ : CascadeMux
    port map (
            O => \N__28536\,
            I => \N__28530\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28527\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28524\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__28527\,
            I => \N__28521\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28518\
        );

    \I__4979\ : Sp12to4
    port map (
            O => \N__28521\,
            I => \N__28515\
        );

    \I__4978\ : Span4Mux_v
    port map (
            O => \N__28518\,
            I => \N__28512\
        );

    \I__4977\ : Odrv12
    port map (
            O => \N__28515\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__28512\,
            I => \current_shift_inst.control_inputZ0Z_21\
        );

    \I__4975\ : InMux
    port map (
            O => \N__28507\,
            I => \current_shift_inst.control_input_1_cry_20\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__28504\,
            I => \N__28501\
        );

    \I__4973\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28498\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28498\,
            I => \N__28495\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__28495\,
            I => \current_shift_inst.control_input_1_axb_6\
        );

    \I__4970\ : CascadeMux
    port map (
            O => \N__28492\,
            I => \N__28489\
        );

    \I__4969\ : InMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__28486\,
            I => \N__28482\
        );

    \I__4967\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28479\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__28482\,
            I => \N__28476\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28473\
        );

    \I__4964\ : Span4Mux_h
    port map (
            O => \N__28476\,
            I => \N__28470\
        );

    \I__4963\ : Odrv12
    port map (
            O => \N__28473\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__4962\ : Odrv4
    port map (
            O => \N__28470\,
            I => \current_shift_inst.control_inputZ0Z_6\
        );

    \I__4961\ : InMux
    port map (
            O => \N__28465\,
            I => \current_shift_inst.control_input_1_cry_5\
        );

    \I__4960\ : CascadeMux
    port map (
            O => \N__28462\,
            I => \N__28459\
        );

    \I__4959\ : InMux
    port map (
            O => \N__28459\,
            I => \N__28456\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__28456\,
            I => \N__28453\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__28453\,
            I => \current_shift_inst.control_input_1_axb_7\
        );

    \I__4956\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28446\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__28449\,
            I => \N__28443\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28440\
        );

    \I__4953\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28437\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__28440\,
            I => \N__28434\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28431\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__28434\,
            I => \N__28428\
        );

    \I__4949\ : Span4Mux_v
    port map (
            O => \N__28431\,
            I => \N__28425\
        );

    \I__4948\ : Odrv4
    port map (
            O => \N__28428\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__28425\,
            I => \current_shift_inst.control_inputZ0Z_7\
        );

    \I__4946\ : InMux
    port map (
            O => \N__28420\,
            I => \current_shift_inst.control_input_1_cry_6\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__28417\,
            I => \N__28414\
        );

    \I__4944\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28411\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__28411\,
            I => \current_shift_inst.control_input_1_axb_8\
        );

    \I__4942\ : CascadeMux
    port map (
            O => \N__28408\,
            I => \N__28404\
        );

    \I__4941\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28401\
        );

    \I__4940\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28398\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__28401\,
            I => \N__28395\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__28398\,
            I => \N__28392\
        );

    \I__4937\ : Span12Mux_v
    port map (
            O => \N__28395\,
            I => \N__28389\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__28392\,
            I => \N__28386\
        );

    \I__4935\ : Odrv12
    port map (
            O => \N__28389\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__28386\,
            I => \current_shift_inst.control_inputZ0Z_8\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28381\,
            I => \bfn_11_21_0_\
        );

    \I__4932\ : InMux
    port map (
            O => \N__28378\,
            I => \N__28375\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__28375\,
            I => \N__28372\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__28372\,
            I => \current_shift_inst.control_input_1_axb_9\
        );

    \I__4929\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28365\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__28368\,
            I => \N__28362\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__28365\,
            I => \N__28359\
        );

    \I__4926\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28356\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__28359\,
            I => \N__28351\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__28356\,
            I => \N__28351\
        );

    \I__4923\ : Span4Mux_h
    port map (
            O => \N__28351\,
            I => \N__28348\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__28348\,
            I => \current_shift_inst.control_inputZ0Z_9\
        );

    \I__4921\ : InMux
    port map (
            O => \N__28345\,
            I => \current_shift_inst.control_input_1_cry_8\
        );

    \I__4920\ : InMux
    port map (
            O => \N__28342\,
            I => \N__28339\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__28336\,
            I => \current_shift_inst.control_input_1_axb_10\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__28333\,
            I => \N__28329\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28326\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28323\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__28326\,
            I => \N__28320\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__28323\,
            I => \N__28317\
        );

    \I__4912\ : Span12Mux_s11_h
    port map (
            O => \N__28320\,
            I => \N__28314\
        );

    \I__4911\ : Span4Mux_h
    port map (
            O => \N__28317\,
            I => \N__28311\
        );

    \I__4910\ : Odrv12
    port map (
            O => \N__28314\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__28311\,
            I => \current_shift_inst.control_inputZ0Z_10\
        );

    \I__4908\ : InMux
    port map (
            O => \N__28306\,
            I => \current_shift_inst.control_input_1_cry_9\
        );

    \I__4907\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28300\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__28297\,
            I => \current_shift_inst.control_input_1_axb_11\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__28294\,
            I => \N__28290\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28287\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28290\,
            I => \N__28284\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__28287\,
            I => \N__28281\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__28284\,
            I => \N__28278\
        );

    \I__4899\ : Span12Mux_s11_h
    port map (
            O => \N__28281\,
            I => \N__28275\
        );

    \I__4898\ : Span4Mux_v
    port map (
            O => \N__28278\,
            I => \N__28272\
        );

    \I__4897\ : Odrv12
    port map (
            O => \N__28275\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__28272\,
            I => \current_shift_inst.control_inputZ0Z_11\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28267\,
            I => \current_shift_inst.control_input_1_cry_10\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28261\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__28261\,
            I => \N__28258\
        );

    \I__4892\ : Odrv4
    port map (
            O => \N__28258\,
            I => \current_shift_inst.control_input_1_axb_12\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__28255\,
            I => \N__28251\
        );

    \I__4890\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28248\
        );

    \I__4889\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28245\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__28248\,
            I => \N__28240\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__28245\,
            I => \N__28240\
        );

    \I__4886\ : Span4Mux_v
    port map (
            O => \N__28240\,
            I => \N__28237\
        );

    \I__4885\ : Odrv4
    port map (
            O => \N__28237\,
            I => \current_shift_inst.control_inputZ0Z_12\
        );

    \I__4884\ : InMux
    port map (
            O => \N__28234\,
            I => \current_shift_inst.control_input_1_cry_11\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28228\,
            I => \N__28225\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__4880\ : Odrv4
    port map (
            O => \N__28222\,
            I => \current_shift_inst.control_input_1_axb_13\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__28219\,
            I => \N__28216\
        );

    \I__4878\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28209\
        );

    \I__4876\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28206\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__28209\,
            I => \N__28203\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__28206\,
            I => \N__28200\
        );

    \I__4873\ : Span4Mux_h
    port map (
            O => \N__28203\,
            I => \N__28197\
        );

    \I__4872\ : Odrv12
    port map (
            O => \N__28200\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__4871\ : Odrv4
    port map (
            O => \N__28197\,
            I => \current_shift_inst.control_inputZ0Z_13\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28192\,
            I => \current_shift_inst.control_input_1_cry_12\
        );

    \I__4869\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28186\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28186\,
            I => \current_shift_inst.control_input_1_axb_0\
        );

    \I__4867\ : InMux
    port map (
            O => \N__28183\,
            I => \N__28180\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__28180\,
            I => \N__28176\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__28179\,
            I => \N__28173\
        );

    \I__4864\ : Span4Mux_v
    port map (
            O => \N__28176\,
            I => \N__28170\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28167\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__28170\,
            I => \N__28162\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28167\,
            I => \N__28162\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__28162\,
            I => \N__28159\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__28159\,
            I => \current_shift_inst.control_inputZ0Z_0\
        );

    \I__4858\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28153\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28153\,
            I => \N__28150\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__28150\,
            I => \current_shift_inst.control_input_1_axb_1\
        );

    \I__4855\ : InMux
    port map (
            O => \N__28147\,
            I => \N__28143\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \N__28140\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28143\,
            I => \N__28137\
        );

    \I__4852\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28134\
        );

    \I__4851\ : Span4Mux_h
    port map (
            O => \N__28137\,
            I => \N__28131\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__28134\,
            I => \N__28128\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__28131\,
            I => \N__28125\
        );

    \I__4848\ : Span4Mux_h
    port map (
            O => \N__28128\,
            I => \N__28122\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__28125\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__28122\,
            I => \current_shift_inst.control_inputZ0Z_1\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28117\,
            I => \current_shift_inst.control_input_1_cry_0\
        );

    \I__4844\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28111\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__28111\,
            I => \N__28108\
        );

    \I__4842\ : Odrv4
    port map (
            O => \N__28108\,
            I => \current_shift_inst.control_input_1_axb_2\
        );

    \I__4841\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28102\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28102\,
            I => \N__28098\
        );

    \I__4839\ : CascadeMux
    port map (
            O => \N__28101\,
            I => \N__28095\
        );

    \I__4838\ : Span4Mux_s3_h
    port map (
            O => \N__28098\,
            I => \N__28092\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28089\
        );

    \I__4836\ : Span4Mux_h
    port map (
            O => \N__28092\,
            I => \N__28086\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__28089\,
            I => \N__28083\
        );

    \I__4834\ : Span4Mux_h
    port map (
            O => \N__28086\,
            I => \N__28080\
        );

    \I__4833\ : Span4Mux_v
    port map (
            O => \N__28083\,
            I => \N__28077\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__28080\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__28077\,
            I => \current_shift_inst.control_inputZ0Z_2\
        );

    \I__4830\ : InMux
    port map (
            O => \N__28072\,
            I => \current_shift_inst.control_input_1_cry_1\
        );

    \I__4829\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28066\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28063\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__28063\,
            I => \current_shift_inst.control_input_1_axb_3\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28057\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28053\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__28056\,
            I => \N__28050\
        );

    \I__4823\ : Span4Mux_h
    port map (
            O => \N__28053\,
            I => \N__28047\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28044\
        );

    \I__4821\ : Span4Mux_h
    port map (
            O => \N__28047\,
            I => \N__28041\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__28044\,
            I => \N__28038\
        );

    \I__4819\ : Sp12to4
    port map (
            O => \N__28041\,
            I => \N__28035\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__28038\,
            I => \N__28032\
        );

    \I__4817\ : Odrv12
    port map (
            O => \N__28035\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__28032\,
            I => \current_shift_inst.control_inputZ0Z_3\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28027\,
            I => \current_shift_inst.control_input_1_cry_2\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__28024\,
            I => \N__28021\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28021\,
            I => \N__28018\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__28018\,
            I => \N__28015\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__28015\,
            I => \current_shift_inst.control_input_1_axb_4\
        );

    \I__4810\ : InMux
    port map (
            O => \N__28012\,
            I => \N__28008\
        );

    \I__4809\ : CascadeMux
    port map (
            O => \N__28011\,
            I => \N__28005\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__28008\,
            I => \N__28002\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28005\,
            I => \N__27999\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__28002\,
            I => \N__27996\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__27999\,
            I => \N__27993\
        );

    \I__4804\ : Span4Mux_h
    port map (
            O => \N__27996\,
            I => \N__27990\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__27993\,
            I => \N__27987\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__27990\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__27987\,
            I => \current_shift_inst.control_inputZ0Z_4\
        );

    \I__4800\ : InMux
    port map (
            O => \N__27982\,
            I => \current_shift_inst.control_input_1_cry_3\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__27979\,
            I => \N__27976\
        );

    \I__4798\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27973\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__27973\,
            I => \N__27970\
        );

    \I__4796\ : Odrv4
    port map (
            O => \N__27970\,
            I => \current_shift_inst.control_input_1_axb_5\
        );

    \I__4795\ : InMux
    port map (
            O => \N__27967\,
            I => \N__27964\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__27964\,
            I => \N__27960\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__27963\,
            I => \N__27957\
        );

    \I__4792\ : Span4Mux_h
    port map (
            O => \N__27960\,
            I => \N__27954\
        );

    \I__4791\ : InMux
    port map (
            O => \N__27957\,
            I => \N__27951\
        );

    \I__4790\ : Span4Mux_v
    port map (
            O => \N__27954\,
            I => \N__27946\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__27951\,
            I => \N__27946\
        );

    \I__4788\ : Span4Mux_v
    port map (
            O => \N__27946\,
            I => \N__27943\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__27943\,
            I => \current_shift_inst.control_inputZ0Z_5\
        );

    \I__4786\ : InMux
    port map (
            O => \N__27940\,
            I => \current_shift_inst.control_input_1_cry_4\
        );

    \I__4785\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27931\
        );

    \I__4784\ : InMux
    port map (
            O => \N__27936\,
            I => \N__27931\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27924\
        );

    \I__4782\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27921\
        );

    \I__4781\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27916\
        );

    \I__4780\ : InMux
    port map (
            O => \N__27928\,
            I => \N__27916\
        );

    \I__4779\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27912\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__27924\,
            I => \N__27909\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__27921\,
            I => \N__27906\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__27916\,
            I => \N__27903\
        );

    \I__4775\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27900\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__27912\,
            I => \N__27897\
        );

    \I__4773\ : Span4Mux_h
    port map (
            O => \N__27909\,
            I => \N__27894\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__27906\,
            I => \N__27891\
        );

    \I__4771\ : Span4Mux_h
    port map (
            O => \N__27903\,
            I => \N__27888\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__27900\,
            I => \N__27885\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__27897\,
            I => \N__27882\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__27894\,
            I => \N__27879\
        );

    \I__4767\ : Span4Mux_v
    port map (
            O => \N__27891\,
            I => \N__27876\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__27888\,
            I => \N__27873\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__27885\,
            I => \N__27868\
        );

    \I__4764\ : Span4Mux_v
    port map (
            O => \N__27882\,
            I => \N__27868\
        );

    \I__4763\ : Odrv4
    port map (
            O => \N__27879\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__27876\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__4761\ : Odrv4
    port map (
            O => \N__27873\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__27868\,
            I => \current_shift_inst.S1_riseZ0\
        );

    \I__4759\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27856\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__27856\,
            I => \current_shift_inst.S1_syncZ0Z0\
        );

    \I__4757\ : InMux
    port map (
            O => \N__27853\,
            I => \N__27850\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__27850\,
            I => \phase_controller_inst1.start_timer_tr_0_sqmuxa\
        );

    \I__4755\ : InMux
    port map (
            O => \N__27847\,
            I => \N__27841\
        );

    \I__4754\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27841\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__27841\,
            I => \current_shift_inst.S1_syncZ0Z1\
        );

    \I__4752\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__27835\,
            I => \current_shift_inst.S1_sync_prevZ0\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__4749\ : InMux
    port map (
            O => \N__27829\,
            I => \N__27826\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__27826\,
            I => \N__27823\
        );

    \I__4747\ : Span4Mux_v
    port map (
            O => \N__27823\,
            I => \N__27820\
        );

    \I__4746\ : Odrv4
    port map (
            O => \N__27820\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\
        );

    \I__4745\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27814\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27811\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__4742\ : Sp12to4
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__4741\ : Odrv12
    port map (
            O => \N__27805\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__27802\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\
        );

    \I__4739\ : InMux
    port map (
            O => \N__27799\,
            I => \N__27796\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__27796\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\
        );

    \I__4737\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27788\
        );

    \I__4736\ : InMux
    port map (
            O => \N__27792\,
            I => \N__27785\
        );

    \I__4735\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27782\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__27788\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__27785\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__27782\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4731\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27770\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27767\
        );

    \I__4729\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27764\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__27770\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27767\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__27764\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4725\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27752\
        );

    \I__4724\ : InMux
    port map (
            O => \N__27756\,
            I => \N__27749\
        );

    \I__4723\ : InMux
    port map (
            O => \N__27755\,
            I => \N__27746\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__27752\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27749\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__27746\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4719\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27734\
        );

    \I__4718\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27731\
        );

    \I__4717\ : InMux
    port map (
            O => \N__27737\,
            I => \N__27728\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__27734\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__27731\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__27728\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4713\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27716\
        );

    \I__4712\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27713\
        );

    \I__4711\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27710\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__27716\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__27713\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__27710\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4707\ : CascadeMux
    port map (
            O => \N__27703\,
            I => \pwm_generator_inst.un1_counterlto9_2_cascade_\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27682\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27682\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27698\,
            I => \N__27682\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27697\,
            I => \N__27682\
        );

    \I__4702\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27677\
        );

    \I__4701\ : InMux
    port map (
            O => \N__27695\,
            I => \N__27677\
        );

    \I__4700\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27668\
        );

    \I__4699\ : InMux
    port map (
            O => \N__27693\,
            I => \N__27668\
        );

    \I__4698\ : InMux
    port map (
            O => \N__27692\,
            I => \N__27668\
        );

    \I__4697\ : InMux
    port map (
            O => \N__27691\,
            I => \N__27668\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__27682\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__27677\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__27668\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27661\,
            I => \N__27656\
        );

    \I__4692\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27653\
        );

    \I__4691\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27650\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__27656\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__27653\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__27650\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27638\
        );

    \I__4686\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27635\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27641\,
            I => \N__27632\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__27638\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__27635\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__27632\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27620\
        );

    \I__4680\ : InMux
    port map (
            O => \N__27624\,
            I => \N__27617\
        );

    \I__4679\ : InMux
    port map (
            O => \N__27623\,
            I => \N__27614\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__27620\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__27617\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__27614\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4675\ : InMux
    port map (
            O => \N__27607\,
            I => \N__27602\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27599\
        );

    \I__4673\ : InMux
    port map (
            O => \N__27605\,
            I => \N__27596\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__27602\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__27599\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__27596\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__27589\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__4668\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27581\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27585\,
            I => \N__27578\
        );

    \I__4666\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27575\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__27581\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__27578\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__27575\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4662\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27565\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__27565\,
            I => \pwm_generator_inst.un1_counterlt9\
        );

    \I__4660\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27559\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27556\
        );

    \I__4658\ : Odrv12
    port map (
            O => \N__27556\,
            I => \il_min_comp1_D1\
        );

    \I__4657\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27549\
        );

    \I__4656\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27546\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__27549\,
            I => \N__27543\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__27546\,
            I => \N__27540\
        );

    \I__4653\ : Span4Mux_h
    port map (
            O => \N__27543\,
            I => \N__27537\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__27540\,
            I => \phase_controller_inst1.N_231\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__27537\,
            I => \phase_controller_inst1.N_231\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27529\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__27529\,
            I => \N__27523\
        );

    \I__4648\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27520\
        );

    \I__4647\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27517\
        );

    \I__4646\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27514\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__27523\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__27520\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__27517\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__27514\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__4641\ : InMux
    port map (
            O => \N__27505\,
            I => \N__27502\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__27502\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\
        );

    \I__4639\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27496\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__27496\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__27493\,
            I => \N__27490\
        );

    \I__4636\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27487\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__27487\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__27484\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_\
        );

    \I__4633\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27478\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__27478\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\
        );

    \I__4631\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27472\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__27472\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\
        );

    \I__4629\ : InMux
    port map (
            O => \N__27469\,
            I => \N__27463\
        );

    \I__4628\ : InMux
    port map (
            O => \N__27468\,
            I => \N__27463\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__27463\,
            I => \N__27460\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__27460\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\
        );

    \I__4625\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27454\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27449\
        );

    \I__4623\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27444\
        );

    \I__4622\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27444\
        );

    \I__4621\ : Span4Mux_h
    port map (
            O => \N__27449\,
            I => \N__27441\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__27444\,
            I => \N__27438\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__27441\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__27438\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\
        );

    \I__4617\ : InMux
    port map (
            O => \N__27433\,
            I => \N__27430\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__27430\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\
        );

    \I__4615\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27424\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__27424\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__4612\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27415\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__27415\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__27412\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_\
        );

    \I__4609\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27406\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__27406\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\
        );

    \I__4607\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27400\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__27400\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__27397\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27394\,
            I => \N__27391\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__27391\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\
        );

    \I__4602\ : CascadeMux
    port map (
            O => \N__27388\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\
        );

    \I__4601\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27382\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__27382\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\
        );

    \I__4599\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27373\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27378\,
            I => \N__27373\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27373\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1\
        );

    \I__4596\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__27367\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14\
        );

    \I__4594\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__27361\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\
        );

    \I__4592\ : CascadeMux
    port map (
            O => \N__27358\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0_cascade_\
        );

    \I__4591\ : InMux
    port map (
            O => \N__27355\,
            I => \current_shift_inst.un38_control_input_0_cry_28\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27352\,
            I => \current_shift_inst.un38_control_input_0_cry_29\
        );

    \I__4589\ : InMux
    port map (
            O => \N__27349\,
            I => \bfn_10_25_0_\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__27346\,
            I => \N__27338\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__27345\,
            I => \N__27334\
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__27344\,
            I => \N__27330\
        );

    \I__4585\ : InMux
    port map (
            O => \N__27343\,
            I => \N__27327\
        );

    \I__4584\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27312\
        );

    \I__4583\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27312\
        );

    \I__4582\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27312\
        );

    \I__4581\ : InMux
    port map (
            O => \N__27337\,
            I => \N__27312\
        );

    \I__4580\ : InMux
    port map (
            O => \N__27334\,
            I => \N__27312\
        );

    \I__4579\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27312\
        );

    \I__4578\ : InMux
    port map (
            O => \N__27330\,
            I => \N__27312\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27327\,
            I => \N__27309\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__27312\,
            I => \N__27306\
        );

    \I__4575\ : Span4Mux_h
    port map (
            O => \N__27309\,
            I => \N__27303\
        );

    \I__4574\ : Span4Mux_v
    port map (
            O => \N__27306\,
            I => \N__27300\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__27303\,
            I => \N__27297\
        );

    \I__4572\ : Span4Mux_v
    port map (
            O => \N__27300\,
            I => \N__27294\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__27297\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__27294\,
            I => \current_shift_inst.control_inputZ0Z_25\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27286\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__27286\,
            I => \N__27283\
        );

    \I__4567\ : Span4Mux_h
    port map (
            O => \N__27283\,
            I => \N__27280\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__27280\,
            I => \N__27277\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__27277\,
            I => il_max_comp2_c
        );

    \I__4564\ : InMux
    port map (
            O => \N__27274\,
            I => \N__27269\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27266\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27272\,
            I => \N__27263\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__27269\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__27266\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__27263\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4558\ : IoInMux
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__27253\,
            I => \N__27250\
        );

    \I__4556\ : Span4Mux_s1_v
    port map (
            O => \N__27250\,
            I => \N__27247\
        );

    \I__4555\ : Odrv4
    port map (
            O => \N__27247\,
            I => \delay_measurement_inst.delay_hc_timer.N_336_i\
        );

    \I__4554\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27240\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27237\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__27240\,
            I => measured_delay_hc_27
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__27237\,
            I => measured_delay_hc_27
        );

    \I__4550\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27228\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27231\,
            I => \N__27225\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__27228\,
            I => measured_delay_hc_28
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__27225\,
            I => measured_delay_hc_28
        );

    \I__4546\ : InMux
    port map (
            O => \N__27220\,
            I => \N__27217\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__27217\,
            I => \N__27214\
        );

    \I__4544\ : Span12Mux_h
    port map (
            O => \N__27214\,
            I => \N__27211\
        );

    \I__4543\ : Odrv12
    port map (
            O => \N__27211\,
            I => il_min_comp1_c
        );

    \I__4542\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27205\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__27205\,
            I => \N__27202\
        );

    \I__4540\ : Odrv12
    port map (
            O => \N__27202\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__27199\,
            I => \N__27196\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__4536\ : Odrv12
    port map (
            O => \N__27190\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27187\,
            I => \current_shift_inst.un38_control_input_0_cry_20\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27184\,
            I => \N__27181\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__27181\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__27178\,
            I => \N__27175\
        );

    \I__4531\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27172\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__4529\ : Odrv12
    port map (
            O => \N__27169\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27166\,
            I => \current_shift_inst.un38_control_input_0_cry_21\
        );

    \I__4527\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27160\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27157\
        );

    \I__4525\ : Span4Mux_v
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__4524\ : Span4Mux_v
    port map (
            O => \N__27154\,
            I => \N__27151\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__27151\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\
        );

    \I__4522\ : CascadeMux
    port map (
            O => \N__27148\,
            I => \N__27145\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27142\,
            I => \N__27139\
        );

    \I__4519\ : Span4Mux_v
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__4518\ : Span4Mux_v
    port map (
            O => \N__27136\,
            I => \N__27133\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__27133\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\
        );

    \I__4516\ : InMux
    port map (
            O => \N__27130\,
            I => \bfn_10_24_0_\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27127\,
            I => \current_shift_inst.un38_control_input_0_cry_23\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27124\,
            I => \current_shift_inst.un38_control_input_0_cry_24\
        );

    \I__4513\ : InMux
    port map (
            O => \N__27121\,
            I => \current_shift_inst.un38_control_input_0_cry_25\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27118\,
            I => \current_shift_inst.un38_control_input_0_cry_26\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27115\,
            I => \current_shift_inst.un38_control_input_0_cry_27\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__27112\,
            I => \N__27109\
        );

    \I__4509\ : InMux
    port map (
            O => \N__27109\,
            I => \N__27106\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__27106\,
            I => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27103\,
            I => \current_shift_inst.un38_control_input_0_cry_11\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__27100\,
            I => \N__27097\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27094\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__27094\,
            I => \N__27091\
        );

    \I__4503\ : Odrv12
    port map (
            O => \N__27091\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27088\,
            I => \current_shift_inst.un38_control_input_0_cry_12\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27082\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__27082\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\
        );

    \I__4499\ : CascadeMux
    port map (
            O => \N__27079\,
            I => \N__27076\
        );

    \I__4498\ : InMux
    port map (
            O => \N__27076\,
            I => \N__27073\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__27073\,
            I => \N__27070\
        );

    \I__4496\ : Odrv12
    port map (
            O => \N__27070\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27067\,
            I => \current_shift_inst.un38_control_input_0_cry_13\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27058\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27058\,
            I => \N__27055\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__27055\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\
        );

    \I__4490\ : InMux
    port map (
            O => \N__27052\,
            I => \bfn_10_23_0_\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27046\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27043\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__27043\,
            I => \N__27040\
        );

    \I__4486\ : Odrv4
    port map (
            O => \N__27040\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__27037\,
            I => \N__27034\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27031\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27031\,
            I => \N__27028\
        );

    \I__4482\ : Odrv12
    port map (
            O => \N__27028\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27025\,
            I => \current_shift_inst.un38_control_input_0_cry_15\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27022\,
            I => \current_shift_inst.un38_control_input_0_cry_16\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27019\,
            I => \N__27016\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__4477\ : Odrv12
    port map (
            O => \N__27013\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27010\,
            I => \current_shift_inst.un38_control_input_0_cry_17\
        );

    \I__4475\ : InMux
    port map (
            O => \N__27007\,
            I => \N__27004\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__27004\,
            I => \N__27001\
        );

    \I__4473\ : Odrv12
    port map (
            O => \N__27001\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__26998\,
            I => \N__26995\
        );

    \I__4471\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26992\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__26992\,
            I => \N__26989\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__26989\,
            I => \N__26986\
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__26986\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\
        );

    \I__4467\ : InMux
    port map (
            O => \N__26983\,
            I => \current_shift_inst.un38_control_input_0_cry_18\
        );

    \I__4466\ : InMux
    port map (
            O => \N__26980\,
            I => \current_shift_inst.un38_control_input_0_cry_19\
        );

    \I__4465\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26974\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__26971\,
            I => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\
        );

    \I__4462\ : InMux
    port map (
            O => \N__26968\,
            I => \N__26965\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__26965\,
            I => \N__26962\
        );

    \I__4460\ : Odrv12
    port map (
            O => \N__26962\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__26959\,
            I => \N__26956\
        );

    \I__4458\ : InMux
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__4456\ : Odrv4
    port map (
            O => \N__26950\,
            I => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__4454\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26941\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__26941\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\
        );

    \I__4452\ : InMux
    port map (
            O => \N__26938\,
            I => \current_shift_inst.un38_control_input_0_cry_5\
        );

    \I__4451\ : InMux
    port map (
            O => \N__26935\,
            I => \N__26932\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__26932\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__26929\,
            I => \N__26926\
        );

    \I__4448\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26923\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__26923\,
            I => \N__26920\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__26920\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\
        );

    \I__4445\ : InMux
    port map (
            O => \N__26917\,
            I => \bfn_10_22_0_\
        );

    \I__4444\ : CascadeMux
    port map (
            O => \N__26914\,
            I => \N__26911\
        );

    \I__4443\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26908\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__26908\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\
        );

    \I__4441\ : InMux
    port map (
            O => \N__26905\,
            I => \current_shift_inst.un38_control_input_0_cry_7\
        );

    \I__4440\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26899\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__26899\,
            I => \N__26896\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__26896\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\
        );

    \I__4437\ : InMux
    port map (
            O => \N__26893\,
            I => \current_shift_inst.un38_control_input_0_cry_8\
        );

    \I__4436\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26887\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__26887\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__26884\,
            I => \N__26881\
        );

    \I__4433\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26878\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__26878\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\
        );

    \I__4431\ : InMux
    port map (
            O => \N__26875\,
            I => \current_shift_inst.un38_control_input_0_cry_9\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__26872\,
            I => \N__26869\
        );

    \I__4429\ : InMux
    port map (
            O => \N__26869\,
            I => \N__26866\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__26866\,
            I => \N__26863\
        );

    \I__4427\ : Odrv12
    port map (
            O => \N__26863\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\
        );

    \I__4426\ : InMux
    port map (
            O => \N__26860\,
            I => \current_shift_inst.un38_control_input_0_cry_10\
        );

    \I__4425\ : InMux
    port map (
            O => \N__26857\,
            I => \N__26854\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__26854\,
            I => \current_shift_inst.z_i_0_31\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__26851\,
            I => \N__26848\
        );

    \I__4422\ : InMux
    port map (
            O => \N__26848\,
            I => \N__26845\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__26845\,
            I => \N__26842\
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__26842\,
            I => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__26839\,
            I => \N__26836\
        );

    \I__4418\ : InMux
    port map (
            O => \N__26836\,
            I => \N__26833\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__26833\,
            I => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\
        );

    \I__4416\ : CascadeMux
    port map (
            O => \N__26830\,
            I => \N__26827\
        );

    \I__4415\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26824\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__26824\,
            I => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\
        );

    \I__4413\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26816\
        );

    \I__4412\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26813\
        );

    \I__4411\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26810\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__26816\,
            I => \N__26806\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__26813\,
            I => \N__26803\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__26810\,
            I => \N__26800\
        );

    \I__4407\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26797\
        );

    \I__4406\ : Span4Mux_v
    port map (
            O => \N__26806\,
            I => \N__26792\
        );

    \I__4405\ : Span4Mux_v
    port map (
            O => \N__26803\,
            I => \N__26792\
        );

    \I__4404\ : Odrv12
    port map (
            O => \N__26800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__26797\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__26792\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__26785\,
            I => \N__26780\
        );

    \I__4400\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26777\
        );

    \I__4399\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26773\
        );

    \I__4398\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26770\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__26777\,
            I => \N__26767\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26764\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__26773\,
            I => \N__26761\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__26770\,
            I => \N__26758\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__26767\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__26764\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__26761\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4390\ : Odrv12
    port map (
            O => \N__26758\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__26749\,
            I => \N__26746\
        );

    \I__4388\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26743\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__26743\,
            I => \N__26739\
        );

    \I__4386\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26735\
        );

    \I__4385\ : Span4Mux_v
    port map (
            O => \N__26739\,
            I => \N__26732\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__26738\,
            I => \N__26729\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26725\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__26732\,
            I => \N__26722\
        );

    \I__4381\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26719\
        );

    \I__4380\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26716\
        );

    \I__4379\ : Span4Mux_h
    port map (
            O => \N__26725\,
            I => \N__26713\
        );

    \I__4378\ : Odrv4
    port map (
            O => \N__26722\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__26719\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__26716\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4375\ : Odrv4
    port map (
            O => \N__26713\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26701\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__26701\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\
        );

    \I__4372\ : CascadeMux
    port map (
            O => \N__26698\,
            I => \phase_controller_inst1.stoper_tr.N_21_cascade_\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__26695\,
            I => \N__26692\
        );

    \I__4370\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26688\
        );

    \I__4369\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26684\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__26688\,
            I => \N__26681\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26678\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__26684\,
            I => \N__26674\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__26681\,
            I => \N__26671\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__26678\,
            I => \N__26668\
        );

    \I__4363\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26665\
        );

    \I__4362\ : Span4Mux_h
    port map (
            O => \N__26674\,
            I => \N__26662\
        );

    \I__4361\ : Odrv4
    port map (
            O => \N__26671\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4360\ : Odrv4
    port map (
            O => \N__26668\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__26665\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4358\ : Odrv4
    port map (
            O => \N__26662\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__4357\ : InMux
    port map (
            O => \N__26653\,
            I => \N__26650\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__26650\,
            I => \N__26647\
        );

    \I__4355\ : Span4Mux_h
    port map (
            O => \N__26647\,
            I => \N__26643\
        );

    \I__4354\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26638\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__26643\,
            I => \N__26635\
        );

    \I__4352\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26632\
        );

    \I__4351\ : InMux
    port map (
            O => \N__26641\,
            I => \N__26629\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__26638\,
            I => \N__26626\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__26635\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__26632\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__26629\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4346\ : Odrv4
    port map (
            O => \N__26626\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__26617\,
            I => \N__26614\
        );

    \I__4344\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26609\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__26613\,
            I => \N__26606\
        );

    \I__4342\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26603\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__26609\,
            I => \N__26599\
        );

    \I__4340\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26596\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__26603\,
            I => \N__26593\
        );

    \I__4338\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26590\
        );

    \I__4337\ : Span4Mux_h
    port map (
            O => \N__26599\,
            I => \N__26587\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26584\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__26593\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__26590\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__26587\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__26584\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__4331\ : InMux
    port map (
            O => \N__26575\,
            I => \N__26571\
        );

    \I__4330\ : InMux
    port map (
            O => \N__26574\,
            I => \N__26568\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__26571\,
            I => \N__26564\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__26568\,
            I => \N__26560\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26567\,
            I => \N__26557\
        );

    \I__4326\ : Span4Mux_h
    port map (
            O => \N__26564\,
            I => \N__26554\
        );

    \I__4325\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26551\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__26560\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26557\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4322\ : Odrv4
    port map (
            O => \N__26554\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__26551\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__4319\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26536\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__26536\,
            I => \N__26533\
        );

    \I__4317\ : Odrv4
    port map (
            O => \N__26533\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31\
        );

    \I__4316\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26527\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__26527\,
            I => \N__26522\
        );

    \I__4314\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26519\
        );

    \I__4313\ : InMux
    port map (
            O => \N__26525\,
            I => \N__26515\
        );

    \I__4312\ : Span4Mux_v
    port map (
            O => \N__26522\,
            I => \N__26512\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__26519\,
            I => \N__26509\
        );

    \I__4310\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26506\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__26515\,
            I => \N__26503\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__26512\,
            I => \N__26498\
        );

    \I__4307\ : Span4Mux_h
    port map (
            O => \N__26509\,
            I => \N__26498\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__26506\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4305\ : Odrv4
    port map (
            O => \N__26503\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__26498\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__4303\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26486\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26483\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26479\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__26486\,
            I => \N__26476\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__26483\,
            I => \N__26473\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26470\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__26479\,
            I => \N__26467\
        );

    \I__4296\ : Span4Mux_h
    port map (
            O => \N__26476\,
            I => \N__26464\
        );

    \I__4295\ : Odrv12
    port map (
            O => \N__26473\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__26470\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__26467\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4292\ : Odrv4
    port map (
            O => \N__26464\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__26455\,
            I => \N__26450\
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__26454\,
            I => \N__26447\
        );

    \I__4289\ : CascadeMux
    port map (
            O => \N__26453\,
            I => \N__26444\
        );

    \I__4288\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26441\
        );

    \I__4287\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26437\
        );

    \I__4286\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26434\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__26441\,
            I => \N__26431\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__26440\,
            I => \N__26428\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__26437\,
            I => \N__26423\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__26434\,
            I => \N__26423\
        );

    \I__4281\ : Span4Mux_h
    port map (
            O => \N__26431\,
            I => \N__26420\
        );

    \I__4280\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26417\
        );

    \I__4279\ : Span4Mux_v
    port map (
            O => \N__26423\,
            I => \N__26414\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__26420\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__26417\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__26414\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__4275\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26403\
        );

    \I__4274\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26398\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__26403\,
            I => \N__26395\
        );

    \I__4272\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26392\
        );

    \I__4271\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26389\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__26398\,
            I => \N__26386\
        );

    \I__4269\ : Odrv12
    port map (
            O => \N__26395\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__26392\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__26389\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__26386\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__4265\ : InMux
    port map (
            O => \N__26377\,
            I => \N__26372\
        );

    \I__4264\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26369\
        );

    \I__4263\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26366\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26362\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__26369\,
            I => \N__26359\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__26366\,
            I => \N__26356\
        );

    \I__4259\ : InMux
    port map (
            O => \N__26365\,
            I => \N__26353\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__26362\,
            I => \N__26350\
        );

    \I__4257\ : Span4Mux_h
    port map (
            O => \N__26359\,
            I => \N__26347\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__26356\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__26353\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__26350\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4253\ : Odrv4
    port map (
            O => \N__26347\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__4252\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26333\
        );

    \I__4251\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26330\
        );

    \I__4250\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26326\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__26333\,
            I => \N__26323\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__26330\,
            I => \N__26320\
        );

    \I__4247\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26317\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__26326\,
            I => \N__26314\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__26323\,
            I => \N__26311\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__26320\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__26317\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4242\ : Odrv4
    port map (
            O => \N__26314\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__26311\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__26302\,
            I => \N__26298\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__26301\,
            I => \N__26295\
        );

    \I__4238\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26291\
        );

    \I__4237\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26288\
        );

    \I__4236\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26285\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__26291\,
            I => \N__26281\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__26288\,
            I => \N__26278\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__26285\,
            I => \N__26275\
        );

    \I__4232\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26272\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__26281\,
            I => \N__26269\
        );

    \I__4230\ : Span4Mux_h
    port map (
            O => \N__26278\,
            I => \N__26266\
        );

    \I__4229\ : Odrv12
    port map (
            O => \N__26275\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__26272\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__26269\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__26266\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26252\
        );

    \I__4224\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26249\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26245\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__26252\,
            I => \N__26242\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__26249\,
            I => \N__26239\
        );

    \I__4220\ : InMux
    port map (
            O => \N__26248\,
            I => \N__26236\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__26245\,
            I => \N__26233\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__26242\,
            I => \N__26230\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__26239\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4216\ : LocalMux
    port map (
            O => \N__26236\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__26233\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__26230\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26218\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26218\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\
        );

    \I__4211\ : InMux
    port map (
            O => \N__26215\,
            I => \N__26212\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__26212\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__26209\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26200\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26205\,
            I => \N__26200\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__26200\,
            I => \N__26197\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__26197\,
            I => \N__26194\
        );

    \I__4204\ : Odrv4
    port map (
            O => \N__26194\,
            I => \current_shift_inst.PI_CTRL.N_46_21\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__26191\,
            I => \N__26187\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__26190\,
            I => \N__26184\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26181\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26177\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__26181\,
            I => \N__26173\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__26180\,
            I => \N__26170\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26177\,
            I => \N__26167\
        );

    \I__4196\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26164\
        );

    \I__4195\ : Span4Mux_h
    port map (
            O => \N__26173\,
            I => \N__26161\
        );

    \I__4194\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26158\
        );

    \I__4193\ : Span4Mux_h
    port map (
            O => \N__26167\,
            I => \N__26153\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__26164\,
            I => \N__26153\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__26161\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26158\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__26153\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__26146\,
            I => \phase_controller_inst1.N_232_cascade_\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26140\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__26140\,
            I => \N__26135\
        );

    \I__4185\ : InMux
    port map (
            O => \N__26139\,
            I => \N__26132\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26129\
        );

    \I__4183\ : Span4Mux_v
    port map (
            O => \N__26135\,
            I => \N__26126\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__26132\,
            I => \N__26121\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__26129\,
            I => \N__26121\
        );

    \I__4180\ : Span4Mux_v
    port map (
            O => \N__26126\,
            I => \N__26118\
        );

    \I__4179\ : Span12Mux_h
    port map (
            O => \N__26121\,
            I => \N__26115\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__26118\,
            I => \il_max_comp1_D2\
        );

    \I__4177\ : Odrv12
    port map (
            O => \N__26115\,
            I => \il_max_comp1_D2\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26107\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26104\
        );

    \I__4174\ : Odrv4
    port map (
            O => \N__26104\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26101\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__4172\ : InMux
    port map (
            O => \N__26098\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26095\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26092\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26089\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26086\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26083\,
            I => \bfn_10_13_0_\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26080\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__26077\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26071\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26071\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto13\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26068\,
            I => \N__26063\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26060\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26057\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26063\,
            I => measured_delay_hc_19
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__26060\,
            I => measured_delay_hc_19
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__26057\,
            I => measured_delay_hc_19
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__26050\,
            I => \N__26047\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__26044\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26041\,
            I => \bfn_10_12_0_\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26038\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__26035\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_\
        );

    \I__4150\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__26029\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__26026\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30_cascade_\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26020\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__26020\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26017\,
            I => \N__26014\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__26014\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__4143\ : CascadeMux
    port map (
            O => \N__26011\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26008\,
            I => \N__26003\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26007\,
            I => \N__26000\
        );

    \I__4140\ : InMux
    port map (
            O => \N__26006\,
            I => \N__25997\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26003\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26000\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__25997\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__4136\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25985\
        );

    \I__4135\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25982\
        );

    \I__4134\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25979\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__25985\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__25982\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__25979\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__4130\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25966\
        );

    \I__4129\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25963\
        );

    \I__4128\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25960\
        );

    \I__4127\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25957\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__25966\,
            I => \N__25952\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__25963\,
            I => \N__25952\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__25960\,
            I => delay_hc_d2
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__25957\,
            I => delay_hc_d2
        );

    \I__4122\ : Odrv4
    port map (
            O => \N__25952\,
            I => delay_hc_d2
        );

    \I__4121\ : InMux
    port map (
            O => \N__25945\,
            I => \N__25941\
        );

    \I__4120\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25938\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__25941\,
            I => measured_delay_hc_26
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__25938\,
            I => measured_delay_hc_26
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__25933\,
            I => \N__25929\
        );

    \I__4116\ : InMux
    port map (
            O => \N__25932\,
            I => \N__25926\
        );

    \I__4115\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25923\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__25926\,
            I => measured_delay_hc_30
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__25923\,
            I => measured_delay_hc_30
        );

    \I__4112\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25914\
        );

    \I__4111\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25911\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__25914\,
            I => measured_delay_hc_25
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__25911\,
            I => measured_delay_hc_25
        );

    \I__4108\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25902\
        );

    \I__4107\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25899\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__25902\,
            I => measured_delay_hc_23
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__25899\,
            I => measured_delay_hc_23
        );

    \I__4104\ : InMux
    port map (
            O => \N__25894\,
            I => \N__25890\
        );

    \I__4103\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25887\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__25890\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__25887\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__4100\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25878\
        );

    \I__4099\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25875\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__25878\,
            I => measured_delay_hc_24
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__25875\,
            I => measured_delay_hc_24
        );

    \I__4096\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25866\
        );

    \I__4095\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25863\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__25866\,
            I => measured_delay_hc_29
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__25863\,
            I => measured_delay_hc_29
        );

    \I__4092\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25855\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25852\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__25852\,
            I => \current_shift_inst.S3_syncZ0Z0\
        );

    \I__4089\ : InMux
    port map (
            O => \N__25849\,
            I => \N__25843\
        );

    \I__4088\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25843\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__25843\,
            I => \current_shift_inst.S3_syncZ0Z1\
        );

    \I__4086\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__25837\,
            I => \current_shift_inst.S3_sync_prevZ0\
        );

    \I__4084\ : InMux
    port map (
            O => \N__25834\,
            I => \N__25831\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__25831\,
            I => \N__25828\
        );

    \I__4082\ : IoSpan4Mux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__25825\,
            I => il_min_comp2_c
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__25822\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3_cascade_\
        );

    \I__4079\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__25816\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\
        );

    \I__4077\ : InMux
    port map (
            O => \N__25813\,
            I => \N__25809\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__25812\,
            I => \N__25806\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__25809\,
            I => \N__25802\
        );

    \I__4074\ : InMux
    port map (
            O => \N__25806\,
            I => \N__25796\
        );

    \I__4073\ : InMux
    port map (
            O => \N__25805\,
            I => \N__25796\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__25802\,
            I => \N__25790\
        );

    \I__4071\ : InMux
    port map (
            O => \N__25801\,
            I => \N__25787\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25784\
        );

    \I__4069\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25779\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25779\
        );

    \I__4067\ : InMux
    port map (
            O => \N__25793\,
            I => \N__25776\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__25790\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__25787\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__25784\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__25779\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__25776\,
            I => \current_shift_inst.meas_stateZ0Z_0\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__25765\,
            I => \N__25762\
        );

    \I__4060\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25758\
        );

    \I__4059\ : CascadeMux
    port map (
            O => \N__25761\,
            I => \N__25754\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__25758\,
            I => \N__25751\
        );

    \I__4057\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25748\
        );

    \I__4056\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25745\
        );

    \I__4055\ : Odrv12
    port map (
            O => \N__25751\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__25748\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__25745\,
            I => \current_shift_inst.S3_riseZ0\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25735\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25735\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__4050\ : CascadeMux
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__4049\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25726\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25726\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__4047\ : InMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__25720\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__25717\,
            I => \N__25714\
        );

    \I__4044\ : InMux
    port map (
            O => \N__25714\,
            I => \N__25711\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__25711\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__25708\,
            I => \N__25700\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25685\
        );

    \I__4040\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25685\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25685\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25685\
        );

    \I__4037\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25685\
        );

    \I__4036\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25678\
        );

    \I__4035\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25678\
        );

    \I__4034\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25678\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__25697\,
            I => \N__25673\
        );

    \I__4032\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25667\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__25685\,
            I => \N__25662\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__25678\,
            I => \N__25662\
        );

    \I__4029\ : InMux
    port map (
            O => \N__25677\,
            I => \N__25659\
        );

    \I__4028\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25646\
        );

    \I__4027\ : InMux
    port map (
            O => \N__25673\,
            I => \N__25637\
        );

    \I__4026\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25637\
        );

    \I__4025\ : InMux
    port map (
            O => \N__25671\,
            I => \N__25637\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25637\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__25667\,
            I => \N__25634\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__25662\,
            I => \N__25631\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25659\,
            I => \N__25628\
        );

    \I__4020\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25623\
        );

    \I__4019\ : InMux
    port map (
            O => \N__25657\,
            I => \N__25623\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__25656\,
            I => \N__25618\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__25655\,
            I => \N__25615\
        );

    \I__4016\ : InMux
    port map (
            O => \N__25654\,
            I => \N__25607\
        );

    \I__4015\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25607\
        );

    \I__4014\ : InMux
    port map (
            O => \N__25652\,
            I => \N__25607\
        );

    \I__4013\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25600\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25600\
        );

    \I__4011\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25600\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__25646\,
            I => \N__25595\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__25637\,
            I => \N__25595\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__25634\,
            I => \N__25586\
        );

    \I__4007\ : Span4Mux_h
    port map (
            O => \N__25631\,
            I => \N__25586\
        );

    \I__4006\ : Span4Mux_v
    port map (
            O => \N__25628\,
            I => \N__25586\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25586\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25575\
        );

    \I__4003\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25575\
        );

    \I__4002\ : InMux
    port map (
            O => \N__25618\,
            I => \N__25575\
        );

    \I__4001\ : InMux
    port map (
            O => \N__25615\,
            I => \N__25575\
        );

    \I__4000\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25575\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__25607\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__25600\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3997\ : Odrv4
    port map (
            O => \N__25595\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__25586\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__25575\,
            I => \current_shift_inst.PI_CTRL.N_75\
        );

    \I__3994\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25561\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__25561\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__25558\,
            I => \N__25555\
        );

    \I__3991\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25541\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__25554\,
            I => \N__25538\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__25553\,
            I => \N__25535\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__25552\,
            I => \N__25532\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__25551\,
            I => \N__25529\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__25550\,
            I => \N__25523\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__25549\,
            I => \N__25517\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__25548\,
            I => \N__25514\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__25547\,
            I => \N__25511\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__25546\,
            I => \N__25506\
        );

    \I__3981\ : CascadeMux
    port map (
            O => \N__25545\,
            I => \N__25503\
        );

    \I__3980\ : CascadeMux
    port map (
            O => \N__25544\,
            I => \N__25500\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25496\
        );

    \I__3978\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25493\
        );

    \I__3977\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25482\
        );

    \I__3976\ : InMux
    port map (
            O => \N__25532\,
            I => \N__25482\
        );

    \I__3975\ : InMux
    port map (
            O => \N__25529\,
            I => \N__25482\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25482\
        );

    \I__3973\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25482\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__25526\,
            I => \N__25479\
        );

    \I__3971\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25470\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__25522\,
            I => \N__25467\
        );

    \I__3969\ : CascadeMux
    port map (
            O => \N__25521\,
            I => \N__25463\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25460\
        );

    \I__3967\ : InMux
    port map (
            O => \N__25517\,
            I => \N__25449\
        );

    \I__3966\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25449\
        );

    \I__3965\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25449\
        );

    \I__3964\ : InMux
    port map (
            O => \N__25510\,
            I => \N__25449\
        );

    \I__3963\ : InMux
    port map (
            O => \N__25509\,
            I => \N__25449\
        );

    \I__3962\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25440\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25440\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25500\,
            I => \N__25440\
        );

    \I__3959\ : InMux
    port map (
            O => \N__25499\,
            I => \N__25440\
        );

    \I__3958\ : Span4Mux_h
    port map (
            O => \N__25496\,
            I => \N__25433\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__25493\,
            I => \N__25433\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__25482\,
            I => \N__25433\
        );

    \I__3955\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25428\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25428\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__25477\,
            I => \N__25425\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__25476\,
            I => \N__25422\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__25475\,
            I => \N__25418\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__25474\,
            I => \N__25414\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__25473\,
            I => \N__25411\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__25470\,
            I => \N__25407\
        );

    \I__3947\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25402\
        );

    \I__3946\ : InMux
    port map (
            O => \N__25466\,
            I => \N__25402\
        );

    \I__3945\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25398\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__25460\,
            I => \N__25395\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__25449\,
            I => \N__25386\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__25440\,
            I => \N__25386\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__25433\,
            I => \N__25386\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__25428\,
            I => \N__25386\
        );

    \I__3939\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25379\
        );

    \I__3938\ : InMux
    port map (
            O => \N__25422\,
            I => \N__25379\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25379\
        );

    \I__3936\ : InMux
    port map (
            O => \N__25418\,
            I => \N__25374\
        );

    \I__3935\ : InMux
    port map (
            O => \N__25417\,
            I => \N__25374\
        );

    \I__3934\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25367\
        );

    \I__3933\ : InMux
    port map (
            O => \N__25411\,
            I => \N__25367\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25367\
        );

    \I__3931\ : Span4Mux_h
    port map (
            O => \N__25407\,
            I => \N__25364\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25402\,
            I => \N__25361\
        );

    \I__3929\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25358\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__25398\,
            I => \N__25351\
        );

    \I__3927\ : Span4Mux_h
    port map (
            O => \N__25395\,
            I => \N__25351\
        );

    \I__3926\ : Span4Mux_v
    port map (
            O => \N__25386\,
            I => \N__25351\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__25379\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__25374\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__25367\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__25364\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3921\ : Odrv12
    port map (
            O => \N__25361\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__25358\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__25351\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3918\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25318\
        );

    \I__3917\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25307\
        );

    \I__3916\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25307\
        );

    \I__3915\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25307\
        );

    \I__3914\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25307\
        );

    \I__3913\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25307\
        );

    \I__3912\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25300\
        );

    \I__3911\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25300\
        );

    \I__3910\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25300\
        );

    \I__3909\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25295\
        );

    \I__3908\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25295\
        );

    \I__3907\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25286\
        );

    \I__3906\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25277\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25277\
        );

    \I__3904\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25277\
        );

    \I__3903\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25277\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__25318\,
            I => \N__25274\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__25307\,
            I => \N__25267\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25300\,
            I => \N__25267\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__25295\,
            I => \N__25267\
        );

    \I__3898\ : InMux
    port map (
            O => \N__25294\,
            I => \N__25264\
        );

    \I__3897\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25253\
        );

    \I__3896\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25253\
        );

    \I__3895\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25253\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25253\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25253\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25242\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25277\,
            I => \N__25242\
        );

    \I__3890\ : Span4Mux_v
    port map (
            O => \N__25274\,
            I => \N__25235\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__25267\,
            I => \N__25235\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__25264\,
            I => \N__25235\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25232\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25252\,
            I => \N__25219\
        );

    \I__3885\ : InMux
    port map (
            O => \N__25251\,
            I => \N__25219\
        );

    \I__3884\ : InMux
    port map (
            O => \N__25250\,
            I => \N__25219\
        );

    \I__3883\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25219\
        );

    \I__3882\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25219\
        );

    \I__3881\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25219\
        );

    \I__3880\ : Odrv12
    port map (
            O => \N__25242\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__25235\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__25232\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25219\,
            I => \current_shift_inst.PI_CTRL.N_76\
        );

    \I__3876\ : CEMux
    port map (
            O => \N__25210\,
            I => \N__25204\
        );

    \I__3875\ : CEMux
    port map (
            O => \N__25209\,
            I => \N__25201\
        );

    \I__3874\ : CEMux
    port map (
            O => \N__25208\,
            I => \N__25198\
        );

    \I__3873\ : CEMux
    port map (
            O => \N__25207\,
            I => \N__25191\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25204\,
            I => \N__25188\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25183\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__25198\,
            I => \N__25183\
        );

    \I__3869\ : CEMux
    port map (
            O => \N__25197\,
            I => \N__25180\
        );

    \I__3868\ : CEMux
    port map (
            O => \N__25196\,
            I => \N__25175\
        );

    \I__3867\ : CEMux
    port map (
            O => \N__25195\,
            I => \N__25169\
        );

    \I__3866\ : CEMux
    port map (
            O => \N__25194\,
            I => \N__25166\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25191\,
            I => \N__25163\
        );

    \I__3864\ : Span4Mux_h
    port map (
            O => \N__25188\,
            I => \N__25156\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__25183\,
            I => \N__25156\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25180\,
            I => \N__25156\
        );

    \I__3861\ : CEMux
    port map (
            O => \N__25179\,
            I => \N__25149\
        );

    \I__3860\ : CEMux
    port map (
            O => \N__25178\,
            I => \N__25146\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__25175\,
            I => \N__25142\
        );

    \I__3858\ : CEMux
    port map (
            O => \N__25174\,
            I => \N__25139\
        );

    \I__3857\ : CEMux
    port map (
            O => \N__25173\,
            I => \N__25136\
        );

    \I__3856\ : CEMux
    port map (
            O => \N__25172\,
            I => \N__25129\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25124\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25166\,
            I => \N__25124\
        );

    \I__3853\ : Span4Mux_h
    port map (
            O => \N__25163\,
            I => \N__25119\
        );

    \I__3852\ : Span4Mux_v
    port map (
            O => \N__25156\,
            I => \N__25119\
        );

    \I__3851\ : CEMux
    port map (
            O => \N__25155\,
            I => \N__25116\
        );

    \I__3850\ : CEMux
    port map (
            O => \N__25154\,
            I => \N__25113\
        );

    \I__3849\ : CEMux
    port map (
            O => \N__25153\,
            I => \N__25110\
        );

    \I__3848\ : CEMux
    port map (
            O => \N__25152\,
            I => \N__25107\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__25149\,
            I => \N__25101\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__25146\,
            I => \N__25101\
        );

    \I__3845\ : CEMux
    port map (
            O => \N__25145\,
            I => \N__25098\
        );

    \I__3844\ : Span4Mux_v
    port map (
            O => \N__25142\,
            I => \N__25091\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__25139\,
            I => \N__25091\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25136\,
            I => \N__25091\
        );

    \I__3841\ : CEMux
    port map (
            O => \N__25135\,
            I => \N__25088\
        );

    \I__3840\ : CEMux
    port map (
            O => \N__25134\,
            I => \N__25085\
        );

    \I__3839\ : CEMux
    port map (
            O => \N__25133\,
            I => \N__25082\
        );

    \I__3838\ : CEMux
    port map (
            O => \N__25132\,
            I => \N__25078\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25074\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__25124\,
            I => \N__25065\
        );

    \I__3835\ : Span4Mux_h
    port map (
            O => \N__25119\,
            I => \N__25065\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__25116\,
            I => \N__25065\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__25113\,
            I => \N__25065\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25110\,
            I => \N__25061\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__25107\,
            I => \N__25058\
        );

    \I__3830\ : CEMux
    port map (
            O => \N__25106\,
            I => \N__25055\
        );

    \I__3829\ : Span4Mux_v
    port map (
            O => \N__25101\,
            I => \N__25049\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25098\,
            I => \N__25049\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__25091\,
            I => \N__25042\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__25088\,
            I => \N__25042\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__25085\,
            I => \N__25042\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__25082\,
            I => \N__25039\
        );

    \I__3823\ : CEMux
    port map (
            O => \N__25081\,
            I => \N__25036\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__25078\,
            I => \N__25033\
        );

    \I__3821\ : CEMux
    port map (
            O => \N__25077\,
            I => \N__25030\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__25074\,
            I => \N__25025\
        );

    \I__3819\ : Span4Mux_v
    port map (
            O => \N__25065\,
            I => \N__25025\
        );

    \I__3818\ : CEMux
    port map (
            O => \N__25064\,
            I => \N__25022\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__25061\,
            I => \N__25015\
        );

    \I__3816\ : Span4Mux_h
    port map (
            O => \N__25058\,
            I => \N__25015\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__25055\,
            I => \N__25015\
        );

    \I__3814\ : CEMux
    port map (
            O => \N__25054\,
            I => \N__25012\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__25049\,
            I => \N__25007\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__25042\,
            I => \N__25007\
        );

    \I__3811\ : Span4Mux_v
    port map (
            O => \N__25039\,
            I => \N__25002\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__25036\,
            I => \N__25002\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__25033\,
            I => \N__24997\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25030\,
            I => \N__24997\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__25025\,
            I => \N__24994\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25022\,
            I => \N__24987\
        );

    \I__3805\ : Sp12to4
    port map (
            O => \N__25015\,
            I => \N__24987\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__24987\
        );

    \I__3803\ : Span4Mux_v
    port map (
            O => \N__25007\,
            I => \N__24980\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__25002\,
            I => \N__24980\
        );

    \I__3801\ : Span4Mux_s2_h
    port map (
            O => \N__24997\,
            I => \N__24980\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__24994\,
            I => \N_717_g\
        );

    \I__3799\ : Odrv12
    port map (
            O => \N__24987\,
            I => \N_717_g\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__24980\,
            I => \N_717_g\
        );

    \I__3797\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24969\
        );

    \I__3796\ : InMux
    port map (
            O => \N__24972\,
            I => \N__24965\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__24969\,
            I => \N__24961\
        );

    \I__3794\ : InMux
    port map (
            O => \N__24968\,
            I => \N__24958\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__24965\,
            I => \N__24955\
        );

    \I__3792\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24952\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__24961\,
            I => \N__24949\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__24958\,
            I => \N__24946\
        );

    \I__3789\ : Odrv12
    port map (
            O => \N__24955\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__24952\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__24949\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__24946\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__3785\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__24934\,
            I => \N__24931\
        );

    \I__3783\ : Span4Mux_v
    port map (
            O => \N__24931\,
            I => \N__24927\
        );

    \I__3782\ : InMux
    port map (
            O => \N__24930\,
            I => \N__24924\
        );

    \I__3781\ : Span4Mux_h
    port map (
            O => \N__24927\,
            I => \N__24919\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24916\
        );

    \I__3779\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24913\
        );

    \I__3778\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24910\
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__24919\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3776\ : Odrv12
    port map (
            O => \N__24916\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__24913\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__24910\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__24901\,
            I => \N__24896\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__24900\,
            I => \N__24893\
        );

    \I__3771\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24890\
        );

    \I__3770\ : InMux
    port map (
            O => \N__24896\,
            I => \N__24887\
        );

    \I__3769\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24884\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__24890\,
            I => \N__24880\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__24887\,
            I => \N__24875\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__24884\,
            I => \N__24875\
        );

    \I__3765\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24872\
        );

    \I__3764\ : Span4Mux_h
    port map (
            O => \N__24880\,
            I => \N__24869\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__24875\,
            I => \N__24866\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__24872\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__24869\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__24866\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__3759\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24853\
        );

    \I__3758\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24853\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__24853\,
            I => \N__24850\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__24850\,
            I => \N__24847\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__24847\,
            I => \current_shift_inst.PI_CTRL.N_46_16\
        );

    \I__3754\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24841\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__24841\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__24838\,
            I => \N__24835\
        );

    \I__3751\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24832\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__24832\,
            I => \N__24829\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__24829\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__3748\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24822\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__24825\,
            I => \N__24818\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__24822\,
            I => \N__24815\
        );

    \I__3745\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24812\
        );

    \I__3744\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24808\
        );

    \I__3743\ : Span4Mux_v
    port map (
            O => \N__24815\,
            I => \N__24803\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__24812\,
            I => \N__24803\
        );

    \I__3741\ : InMux
    port map (
            O => \N__24811\,
            I => \N__24800\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__24808\,
            I => \N__24795\
        );

    \I__3739\ : Span4Mux_h
    port map (
            O => \N__24803\,
            I => \N__24795\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__24800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__24795\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__3736\ : InMux
    port map (
            O => \N__24790\,
            I => \N__24787\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__24787\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__3734\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24781\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__24781\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__3732\ : InMux
    port map (
            O => \N__24778\,
            I => \N__24775\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__24775\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__24772\,
            I => \N__24769\
        );

    \I__3729\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24766\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24766\,
            I => \N__24763\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__24763\,
            I => \N__24760\
        );

    \I__3726\ : Span4Mux_v
    port map (
            O => \N__24760\,
            I => \N__24757\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__24757\,
            I => \pwm_generator_inst.thresholdZ0Z_7\
        );

    \I__3724\ : InMux
    port map (
            O => \N__24754\,
            I => \N__24751\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__24751\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__24748\,
            I => \N__24745\
        );

    \I__3721\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24742\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__3719\ : Span4Mux_h
    port map (
            O => \N__24739\,
            I => \N__24736\
        );

    \I__3718\ : Span4Mux_h
    port map (
            O => \N__24736\,
            I => \N__24733\
        );

    \I__3717\ : Odrv4
    port map (
            O => \N__24733\,
            I => \pwm_generator_inst.thresholdZ0Z_8\
        );

    \I__3716\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24727\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__24727\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__24724\,
            I => \N__24721\
        );

    \I__3713\ : InMux
    port map (
            O => \N__24721\,
            I => \N__24718\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__24718\,
            I => \N__24715\
        );

    \I__3711\ : Span4Mux_v
    port map (
            O => \N__24715\,
            I => \N__24712\
        );

    \I__3710\ : Span4Mux_h
    port map (
            O => \N__24712\,
            I => \N__24709\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__24709\,
            I => \pwm_generator_inst.thresholdZ0Z_9\
        );

    \I__3708\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24703\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__24703\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24700\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__3705\ : IoInMux
    port map (
            O => \N__24697\,
            I => \N__24694\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__3703\ : Span4Mux_s1_v
    port map (
            O => \N__24691\,
            I => \N__24688\
        );

    \I__3702\ : Sp12to4
    port map (
            O => \N__24688\,
            I => \N__24685\
        );

    \I__3701\ : Span12Mux_h
    port map (
            O => \N__24685\,
            I => \N__24682\
        );

    \I__3700\ : Odrv12
    port map (
            O => \N__24682\,
            I => pwm_output_c
        );

    \I__3699\ : CascadeMux
    port map (
            O => \N__24679\,
            I => \N__24676\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24673\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24670\
        );

    \I__3696\ : Odrv12
    port map (
            O => \N__24670\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__3695\ : CascadeMux
    port map (
            O => \N__24667\,
            I => \N__24664\
        );

    \I__3694\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24661\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__24661\,
            I => \N__24658\
        );

    \I__3692\ : Span4Mux_h
    port map (
            O => \N__24658\,
            I => \N__24655\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__24655\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__24652\,
            I => \N__24649\
        );

    \I__3689\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24646\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__24646\,
            I => \N__24643\
        );

    \I__3687\ : Span4Mux_h
    port map (
            O => \N__24643\,
            I => \N__24640\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__24640\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__3685\ : CEMux
    port map (
            O => \N__24637\,
            I => \N__24633\
        );

    \I__3684\ : CEMux
    port map (
            O => \N__24636\,
            I => \N__24630\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24627\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__24630\,
            I => \N__24623\
        );

    \I__3681\ : Span4Mux_v
    port map (
            O => \N__24627\,
            I => \N__24618\
        );

    \I__3680\ : CEMux
    port map (
            O => \N__24626\,
            I => \N__24615\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__24623\,
            I => \N__24612\
        );

    \I__3678\ : CEMux
    port map (
            O => \N__24622\,
            I => \N__24609\
        );

    \I__3677\ : CEMux
    port map (
            O => \N__24621\,
            I => \N__24606\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__24618\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__24615\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__24612\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__24609\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__24606\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__3671\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24591\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24588\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__24591\,
            I => \N__24583\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24580\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24577\
        );

    \I__3666\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24574\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__24583\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__3664\ : Odrv4
    port map (
            O => \N__24580\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__24577\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__24574\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__3660\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__24559\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__3658\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24550\
        );

    \I__3657\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24543\
        );

    \I__3656\ : InMux
    port map (
            O => \N__24554\,
            I => \N__24543\
        );

    \I__3655\ : InMux
    port map (
            O => \N__24553\,
            I => \N__24543\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__24550\,
            I => \N__24536\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__24543\,
            I => \N__24536\
        );

    \I__3652\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24533\
        );

    \I__3651\ : InMux
    port map (
            O => \N__24541\,
            I => \N__24530\
        );

    \I__3650\ : Span4Mux_v
    port map (
            O => \N__24536\,
            I => \N__24525\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__24533\,
            I => \N__24525\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__24530\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__24525\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__24520\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_\
        );

    \I__3645\ : InMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__24514\,
            I => \phase_controller_inst1.stoper_hc.un1_startlt15\
        );

    \I__3643\ : CascadeMux
    port map (
            O => \N__24511\,
            I => \N__24508\
        );

    \I__3642\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24505\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__24505\,
            I => \N__24502\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__24502\,
            I => \N__24499\
        );

    \I__3639\ : Span4Mux_v
    port map (
            O => \N__24499\,
            I => \N__24496\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__24496\,
            I => \pwm_generator_inst.thresholdZ0Z_0\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24490\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24490\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__24487\,
            I => \N__24484\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24481\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__24481\,
            I => \pwm_generator_inst.thresholdZ0Z_1\
        );

    \I__3632\ : InMux
    port map (
            O => \N__24478\,
            I => \N__24475\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__24475\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__24472\,
            I => \N__24469\
        );

    \I__3629\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24466\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24463\
        );

    \I__3627\ : Span4Mux_v
    port map (
            O => \N__24463\,
            I => \N__24460\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__24460\,
            I => \pwm_generator_inst.thresholdZ0Z_2\
        );

    \I__3625\ : InMux
    port map (
            O => \N__24457\,
            I => \N__24454\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24454\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__24451\,
            I => \N__24448\
        );

    \I__3622\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24445\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__24445\,
            I => \pwm_generator_inst.thresholdZ0Z_3\
        );

    \I__3620\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24439\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__24439\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__24436\,
            I => \N__24433\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24430\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24427\
        );

    \I__3615\ : Odrv4
    port map (
            O => \N__24427\,
            I => \pwm_generator_inst.thresholdZ0Z_4\
        );

    \I__3614\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__24421\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__24418\,
            I => \N__24415\
        );

    \I__3611\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24412\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__3609\ : Span4Mux_v
    port map (
            O => \N__24409\,
            I => \N__24406\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__24406\,
            I => \pwm_generator_inst.thresholdZ0Z_5\
        );

    \I__3607\ : InMux
    port map (
            O => \N__24403\,
            I => \N__24400\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__24400\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__24397\,
            I => \N__24394\
        );

    \I__3604\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24391\,
            I => \N__24388\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__24382\,
            I => \pwm_generator_inst.thresholdZ0Z_6\
        );

    \I__3599\ : InMux
    port map (
            O => \N__24379\,
            I => \N__24376\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__24376\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24373\,
            I => \N__24370\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__24370\,
            I => \N__24366\
        );

    \I__3595\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24362\
        );

    \I__3594\ : Span4Mux_v
    port map (
            O => \N__24366\,
            I => \N__24359\
        );

    \I__3593\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24356\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__24362\,
            I => measured_delay_hc_21
        );

    \I__3591\ : Odrv4
    port map (
            O => \N__24359\,
            I => measured_delay_hc_21
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__24356\,
            I => measured_delay_hc_21
        );

    \I__3589\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24344\
        );

    \I__3588\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24341\
        );

    \I__3587\ : InMux
    port map (
            O => \N__24347\,
            I => \N__24338\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__24344\,
            I => measured_delay_hc_20
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__24341\,
            I => measured_delay_hc_20
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__24338\,
            I => measured_delay_hc_20
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__24331\,
            I => \N__24326\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__24330\,
            I => \N__24323\
        );

    \I__3581\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24320\
        );

    \I__3580\ : InMux
    port map (
            O => \N__24326\,
            I => \N__24317\
        );

    \I__3579\ : InMux
    port map (
            O => \N__24323\,
            I => \N__24314\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__24320\,
            I => measured_delay_hc_22
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__24317\,
            I => measured_delay_hc_22
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__24314\,
            I => measured_delay_hc_22
        );

    \I__3575\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24304\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__24304\,
            I => \N__24301\
        );

    \I__3573\ : Span12Mux_h
    port map (
            O => \N__24301\,
            I => \N__24298\
        );

    \I__3572\ : Odrv12
    port map (
            O => \N__24298\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_4\
        );

    \I__3571\ : InMux
    port map (
            O => \N__24295\,
            I => \N__24292\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__24292\,
            I => \N__24289\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__24289\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2\
        );

    \I__3568\ : CascadeMux
    port map (
            O => \N__24286\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24280\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__24280\,
            I => \current_shift_inst.N_199\
        );

    \I__3565\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24274\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__24274\,
            I => \N__24271\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__24271\,
            I => \N__24266\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__24270\,
            I => \N__24263\
        );

    \I__3561\ : InMux
    port map (
            O => \N__24269\,
            I => \N__24259\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__24266\,
            I => \N__24256\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24250\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24250\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24245\
        );

    \I__3556\ : Span4Mux_h
    port map (
            O => \N__24256\,
            I => \N__24245\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24242\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__24250\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__24245\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__24242\,
            I => \current_shift_inst.phase_validZ0\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__24235\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4_cascade_\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24232\,
            I => \N__24229\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__24229\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3\
        );

    \I__3548\ : InMux
    port map (
            O => \N__24226\,
            I => \bfn_8_20_0_\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24223\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24220\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24217\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__3544\ : InMux
    port map (
            O => \N__24214\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__3543\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24208\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__24208\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24205\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__3540\ : InMux
    port map (
            O => \N__24202\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__3539\ : InMux
    port map (
            O => \N__24199\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24193\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24193\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__3536\ : InMux
    port map (
            O => \N__24190\,
            I => \bfn_8_19_0_\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24187\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24184\,
            I => \N__24180\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24176\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__24180\,
            I => \N__24173\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__24179\,
            I => \N__24170\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24164\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__24173\,
            I => \N__24161\
        );

    \I__3528\ : InMux
    port map (
            O => \N__24170\,
            I => \N__24156\
        );

    \I__3527\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24156\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24153\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24167\,
            I => \N__24150\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__24164\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__24161\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__24156\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__24153\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24150\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__3519\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24136\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24136\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24133\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__24130\,
            I => \N__24127\
        );

    \I__3515\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24124\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__24124\,
            I => \N__24121\
        );

    \I__3513\ : Odrv4
    port map (
            O => \N__24121\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24118\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__3511\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24112\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24112\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24109\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24106\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24100\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24100\,
            I => \N__24097\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__24097\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24094\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24088\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__24088\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24085\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24082\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24079\,
            I => \N__24074\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24068\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24068\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24065\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24062\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24059\
        );

    \I__3493\ : Span4Mux_h
    port map (
            O => \N__24065\,
            I => \N__24054\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__24062\,
            I => \N__24054\
        );

    \I__3491\ : Span4Mux_h
    port map (
            O => \N__24059\,
            I => \N__24051\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__24054\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3489\ : Odrv4
    port map (
            O => \N__24051\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24043\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__24043\,
            I => \N__24040\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__24040\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24037\,
            I => \bfn_8_18_0_\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24034\,
            I => \N__24029\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24024\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24032\,
            I => \N__24024\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24021\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__24017\
        );

    \I__3479\ : Span4Mux_h
    port map (
            O => \N__24021\,
            I => \N__24014\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24020\,
            I => \N__24011\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__24017\,
            I => \N__24008\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__24014\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__24011\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__24008\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__23998\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__3471\ : InMux
    port map (
            O => \N__23995\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\
        );

    \I__3470\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23989\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__23989\,
            I => \N__23986\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__23986\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__3467\ : InMux
    port map (
            O => \N__23983\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__3466\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23977\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__23977\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__3464\ : InMux
    port map (
            O => \N__23974\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__3463\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23968\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__23968\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__3461\ : InMux
    port map (
            O => \N__23965\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__3460\ : InMux
    port map (
            O => \N__23962\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__3459\ : InMux
    port map (
            O => \N__23959\,
            I => \N__23956\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__23956\,
            I => \N__23953\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__23953\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__3456\ : InMux
    port map (
            O => \N__23950\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__3455\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23944\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__23944\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__3453\ : InMux
    port map (
            O => \N__23941\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__3452\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23934\
        );

    \I__3451\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23931\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__23934\,
            I => \N__23925\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__23931\,
            I => \N__23925\
        );

    \I__3448\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23922\
        );

    \I__3447\ : Span4Mux_h
    port map (
            O => \N__23925\,
            I => \N__23919\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__23922\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__23919\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_0\
        );

    \I__3444\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23909\
        );

    \I__3443\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23906\
        );

    \I__3442\ : InMux
    port map (
            O => \N__23912\,
            I => \N__23903\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__23909\,
            I => \N__23898\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__23906\,
            I => \N__23898\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__23903\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3438\ : Odrv12
    port map (
            O => \N__23898\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__3437\ : InMux
    port map (
            O => \N__23893\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__23890\,
            I => \N__23886\
        );

    \I__3435\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23882\
        );

    \I__3434\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23879\
        );

    \I__3433\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23876\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23871\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23871\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__23876\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3429\ : Odrv12
    port map (
            O => \N__23871\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__3428\ : InMux
    port map (
            O => \N__23866\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__3427\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__3426\ : InMux
    port map (
            O => \N__23862\,
            I => \N__23850\
        );

    \I__3425\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23850\
        );

    \I__3424\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23850\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__23857\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__23850\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0\
        );

    \I__3421\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23839\
        );

    \I__3420\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23834\
        );

    \I__3419\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23834\
        );

    \I__3418\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23831\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23826\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23826\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__23831\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3414\ : Odrv12
    port map (
            O => \N__23826\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__3413\ : InMux
    port map (
            O => \N__23821\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__23818\,
            I => \N__23813\
        );

    \I__3411\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23808\
        );

    \I__3410\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23808\
        );

    \I__3409\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23805\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23800\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__23805\,
            I => \N__23800\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__23800\,
            I => \N__23797\
        );

    \I__3405\ : Span4Mux_h
    port map (
            O => \N__23797\,
            I => \N__23793\
        );

    \I__3404\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23790\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__23793\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__23790\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23779\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__3398\ : InMux
    port map (
            O => \N__23776\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__3397\ : InMux
    port map (
            O => \N__23773\,
            I => \N__23770\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__23770\,
            I => \N__23766\
        );

    \I__3395\ : InMux
    port map (
            O => \N__23769\,
            I => \N__23761\
        );

    \I__3394\ : Span4Mux_h
    port map (
            O => \N__23766\,
            I => \N__23758\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23753\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23753\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__23761\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__23758\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23753\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__3388\ : InMux
    port map (
            O => \N__23746\,
            I => \N__23743\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__23743\,
            I => \N__23740\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__23740\,
            I => \N__23737\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__23737\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23734\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__3383\ : InMux
    port map (
            O => \N__23731\,
            I => \N__23726\
        );

    \I__3382\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23721\
        );

    \I__3381\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23721\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__23726\,
            I => \N__23715\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__23721\,
            I => \N__23715\
        );

    \I__3378\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23712\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__23715\,
            I => \N__23709\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23712\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__23709\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__3374\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23701\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__23701\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__3372\ : InMux
    port map (
            O => \N__23698\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23691\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__23694\,
            I => \N__23687\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23684\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23679\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23687\,
            I => \N__23679\
        );

    \I__3366\ : Span4Mux_h
    port map (
            O => \N__23684\,
            I => \N__23673\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__23679\,
            I => \N__23673\
        );

    \I__3364\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23670\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__23673\,
            I => \N__23667\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__23670\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__23667\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__3360\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23659\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__23659\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__23656\,
            I => \phase_controller_inst1.N_228_cascade_\
        );

    \I__3357\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__23650\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__3355\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23643\
        );

    \I__3354\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23640\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__23643\,
            I => \N__23637\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__23640\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__23637\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__23632\,
            I => \N__23622\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__23631\,
            I => \N__23618\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__23630\,
            I => \N__23614\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__23629\,
            I => \N__23610\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__23628\,
            I => \N__23606\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \N__23601\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__23626\,
            I => \N__23598\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__23625\,
            I => \N__23594\
        );

    \I__3342\ : InMux
    port map (
            O => \N__23622\,
            I => \N__23579\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23579\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23579\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23579\
        );

    \I__3338\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23579\
        );

    \I__3337\ : InMux
    port map (
            O => \N__23613\,
            I => \N__23579\
        );

    \I__3336\ : InMux
    port map (
            O => \N__23610\,
            I => \N__23579\
        );

    \I__3335\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23560\
        );

    \I__3334\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23560\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23560\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23560\
        );

    \I__3331\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23560\
        );

    \I__3330\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23560\
        );

    \I__3329\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23560\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23594\,
            I => \N__23560\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__23579\,
            I => \N__23557\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__23578\,
            I => \N__23553\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__23577\,
            I => \N__23547\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__23560\,
            I => \N__23544\
        );

    \I__3323\ : Span4Mux_v
    port map (
            O => \N__23557\,
            I => \N__23541\
        );

    \I__3322\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23532\
        );

    \I__3321\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23532\
        );

    \I__3320\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23532\
        );

    \I__3319\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23532\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23524\
        );

    \I__3317\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23524\
        );

    \I__3316\ : Span4Mux_h
    port map (
            O => \N__23544\,
            I => \N__23517\
        );

    \I__3315\ : Span4Mux_h
    port map (
            O => \N__23541\,
            I => \N__23517\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__23532\,
            I => \N__23517\
        );

    \I__3313\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23510\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23510\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23510\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__23524\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__23517\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__23510\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__23503\,
            I => \N__23489\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__23502\,
            I => \N__23485\
        );

    \I__3305\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23466\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23466\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23466\
        );

    \I__3302\ : InMux
    port map (
            O => \N__23498\,
            I => \N__23466\
        );

    \I__3301\ : InMux
    port map (
            O => \N__23497\,
            I => \N__23466\
        );

    \I__3300\ : InMux
    port map (
            O => \N__23496\,
            I => \N__23466\
        );

    \I__3299\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23466\
        );

    \I__3298\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23466\
        );

    \I__3297\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23461\
        );

    \I__3296\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23448\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23448\
        );

    \I__3294\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23448\
        );

    \I__3293\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23448\
        );

    \I__3292\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23448\
        );

    \I__3291\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23448\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__23466\,
            I => \N__23445\
        );

    \I__3289\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23433\
        );

    \I__3288\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23433\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__23461\,
            I => \N__23428\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__23448\,
            I => \N__23428\
        );

    \I__3285\ : Span4Mux_h
    port map (
            O => \N__23445\,
            I => \N__23425\
        );

    \I__3284\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23420\
        );

    \I__3283\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23420\
        );

    \I__3282\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23411\
        );

    \I__3281\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23411\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23411\
        );

    \I__3279\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23411\
        );

    \I__3278\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23408\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__23433\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__23428\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__23425\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__23420\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__23411\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__23408\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__23395\,
            I => \N__23388\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__23394\,
            I => \N__23385\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__23393\,
            I => \N__23382\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__23392\,
            I => \N__23379\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__23391\,
            I => \N__23371\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23356\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23356\
        );

    \I__3264\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23356\
        );

    \I__3263\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23356\
        );

    \I__3262\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23347\
        );

    \I__3261\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23347\
        );

    \I__3260\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23347\
        );

    \I__3259\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23347\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__23374\,
            I => \N__23341\
        );

    \I__3257\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23332\
        );

    \I__3256\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23332\
        );

    \I__3255\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23332\
        );

    \I__3254\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23323\
        );

    \I__3253\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23323\
        );

    \I__3252\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23323\
        );

    \I__3251\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23323\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__23356\,
            I => \N__23318\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__23347\,
            I => \N__23318\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__23346\,
            I => \N__23315\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \N__23311\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__23344\,
            I => \N__23308\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23301\
        );

    \I__3244\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23301\
        );

    \I__3243\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23298\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__23332\,
            I => \N__23293\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__23323\,
            I => \N__23293\
        );

    \I__3240\ : Span4Mux_h
    port map (
            O => \N__23318\,
            I => \N__23290\
        );

    \I__3239\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23285\
        );

    \I__3238\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23285\
        );

    \I__3237\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23278\
        );

    \I__3236\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23278\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23278\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23275\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__23301\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__23298\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3231\ : Odrv12
    port map (
            O => \N__23293\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__23290\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23285\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__23278\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__23275\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3226\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23257\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__23257\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23251\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23247\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23244\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__23247\,
            I => \N__23241\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__23244\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__23241\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23236\,
            I => \N__23233\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__23233\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23226\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23223\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23220\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__23223\,
            I => \N__23217\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__23220\,
            I => \N__23214\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__23217\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__23214\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__23206\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__3207\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23200\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__23200\,
            I => \N__23196\
        );

    \I__3205\ : InMux
    port map (
            O => \N__23199\,
            I => \N__23193\
        );

    \I__3204\ : Span4Mux_h
    port map (
            O => \N__23196\,
            I => \N__23190\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23193\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3202\ : Odrv4
    port map (
            O => \N__23190\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3201\ : InMux
    port map (
            O => \N__23185\,
            I => \N__23182\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__23182\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23173\
        );

    \I__3197\ : Span4Mux_h
    port map (
            O => \N__23173\,
            I => \N__23170\
        );

    \I__3196\ : Span4Mux_h
    port map (
            O => \N__23170\,
            I => \N__23167\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__23167\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_3\
        );

    \I__3194\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23161\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__23161\,
            I => \N__23158\
        );

    \I__3192\ : Span4Mux_h
    port map (
            O => \N__23158\,
            I => \N__23155\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__23155\,
            I => \N__23152\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__23152\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_1\
        );

    \I__3189\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23146\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__23146\,
            I => \N__23143\
        );

    \I__3187\ : Span4Mux_v
    port map (
            O => \N__23143\,
            I => \N__23140\
        );

    \I__3186\ : Span4Mux_h
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__23137\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__23134\,
            I => \N__23131\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23128\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23125\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__23122\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23116\,
            I => \N__23113\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__23113\,
            I => \N__23110\
        );

    \I__3176\ : Span4Mux_v
    port map (
            O => \N__23110\,
            I => \N__23107\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__23107\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23101\,
            I => \N__23098\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23095\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__23092\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__3168\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23083\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__23083\,
            I => \N__23080\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__3164\ : Odrv4
    port map (
            O => \N__23074\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__23071\,
            I => \N__23068\
        );

    \I__3162\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23065\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__23062\
        );

    \I__3160\ : Span4Mux_h
    port map (
            O => \N__23062\,
            I => \N__23059\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__23059\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__3158\ : IoInMux
    port map (
            O => \N__23056\,
            I => \N__23053\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23053\,
            I => \N__23050\
        );

    \I__3156\ : IoSpan4Mux
    port map (
            O => \N__23050\,
            I => \N__23047\
        );

    \I__3155\ : Span4Mux_s2_v
    port map (
            O => \N__23047\,
            I => \N__23044\
        );

    \I__3154\ : Span4Mux_v
    port map (
            O => \N__23044\,
            I => \N__23041\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__23041\,
            I => \current_shift_inst.timer_s1.N_187_i\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23038\,
            I => \N__23035\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__3150\ : Odrv12
    port map (
            O => \N__23032\,
            I => il_max_comp1_c
        );

    \I__3149\ : InMux
    port map (
            O => \N__23029\,
            I => \N__23026\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__3147\ : Odrv12
    port map (
            O => \N__23023\,
            I => \il_max_comp1_D1\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23017\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23014\
        );

    \I__3144\ : Odrv12
    port map (
            O => \N__23014\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_7\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23008\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__3141\ : Odrv12
    port map (
            O => \N__23005\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_2\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__3139\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22996\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__22996\,
            I => \N__22993\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__22993\,
            I => \N__22990\
        );

    \I__3136\ : Span4Mux_h
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__22987\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__22984\,
            I => \N__22981\
        );

    \I__3133\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__22978\,
            I => \N__22975\
        );

    \I__3131\ : Span4Mux_h
    port map (
            O => \N__22975\,
            I => \N__22972\
        );

    \I__3130\ : Odrv4
    port map (
            O => \N__22972\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__22969\,
            I => \N__22966\
        );

    \I__3128\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22963\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22960\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__22957\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__3123\ : InMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__22945\,
            I => \N__22942\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__22942\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__3118\ : InMux
    port map (
            O => \N__22936\,
            I => \N__22933\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__22930\,
            I => \N__22927\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__22927\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__3114\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__22921\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31\
        );

    \I__3112\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__22915\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2\
        );

    \I__3110\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22909\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22905\
        );

    \I__3108\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22902\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__22905\,
            I => \N__22897\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__22902\,
            I => \N__22897\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__22897\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__22894\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_\
        );

    \I__3103\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22885\
        );

    \I__3102\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22885\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__22885\,
            I => \N__22882\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__22882\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__3099\ : InMux
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__22876\,
            I => \N__22872\
        );

    \I__3097\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22869\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__22872\,
            I => \N__22866\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22863\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__22866\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3093\ : Odrv12
    port map (
            O => \N__22863\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3092\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22855\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22852\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__22852\,
            I => \N__22849\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__22849\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__3088\ : InMux
    port map (
            O => \N__22846\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__3087\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22840\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__22840\,
            I => \N__22836\
        );

    \I__3085\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22833\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__22836\,
            I => \N__22828\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__22833\,
            I => \N__22828\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__22828\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__3081\ : InMux
    port map (
            O => \N__22825\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__3080\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22819\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__22819\,
            I => \N__22816\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__22816\,
            I => \N__22813\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__22813\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__3076\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22807\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__22807\,
            I => \N__22804\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__22804\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \current_shift_inst.PI_CTRL.N_47_16_cascade_\
        );

    \I__3072\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22795\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22792\
        );

    \I__3070\ : Odrv12
    port map (
            O => \N__22792\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\
        );

    \I__3069\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22786\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__22786\,
            I => \current_shift_inst.PI_CTRL.N_47_21\
        );

    \I__3067\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__22780\,
            I => \current_shift_inst.PI_CTRL.N_47_16\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__22777\,
            I => \current_shift_inst.PI_CTRL.N_47_21_cascade_\
        );

    \I__3064\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22771\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__22771\,
            I => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\
        );

    \I__3062\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22765\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__22765\,
            I => \N__22761\
        );

    \I__3060\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22758\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__22761\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__22758\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3057\ : InMux
    port map (
            O => \N__22753\,
            I => \N__22750\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__3055\ : Odrv12
    port map (
            O => \N__22747\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__3054\ : InMux
    port map (
            O => \N__22744\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22738\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__22738\,
            I => \N__22734\
        );

    \I__3051\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22731\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__22734\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__22731\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3048\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__22723\,
            I => \N__22720\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__22720\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__3045\ : InMux
    port map (
            O => \N__22717\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22711\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22707\
        );

    \I__3042\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22704\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__22707\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__22704\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3039\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22696\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__22696\,
            I => \N__22693\
        );

    \I__3037\ : Odrv4
    port map (
            O => \N__22693\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__3036\ : InMux
    port map (
            O => \N__22690\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__3035\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22683\
        );

    \I__3034\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22680\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22677\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__22680\,
            I => \N__22674\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__22677\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3030\ : Odrv4
    port map (
            O => \N__22674\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3029\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22666\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__22666\,
            I => \N__22663\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__22663\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__3026\ : InMux
    port map (
            O => \N__22660\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__3025\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22650\
        );

    \I__3023\ : InMux
    port map (
            O => \N__22653\,
            I => \N__22647\
        );

    \I__3022\ : Odrv12
    port map (
            O => \N__22650\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__22647\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3020\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22639\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__22636\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__3017\ : InMux
    port map (
            O => \N__22633\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__3016\ : InMux
    port map (
            O => \N__22630\,
            I => \N__22627\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22624\
        );

    \I__3014\ : Span4Mux_h
    port map (
            O => \N__22624\,
            I => \N__22620\
        );

    \I__3013\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22617\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__22620\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__22617\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3010\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22609\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__22609\,
            I => \N__22606\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__22606\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__3007\ : InMux
    port map (
            O => \N__22603\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__3006\ : InMux
    port map (
            O => \N__22600\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__3005\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22594\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__22594\,
            I => \N__22590\
        );

    \I__3003\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22587\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__22590\,
            I => \N__22584\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__22587\,
            I => \N__22581\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__22584\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2999\ : Odrv12
    port map (
            O => \N__22581\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__2998\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22573\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__22573\,
            I => \N__22570\
        );

    \I__2996\ : Span4Mux_h
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__22567\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__2994\ : InMux
    port map (
            O => \N__22564\,
            I => \bfn_7_15_0_\
        );

    \I__2993\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22558\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__22558\,
            I => \N__22555\
        );

    \I__2991\ : Span4Mux_h
    port map (
            O => \N__22555\,
            I => \N__22551\
        );

    \I__2990\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22548\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__22551\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__22548\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__2987\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__22540\,
            I => \N__22537\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__22534\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__2983\ : InMux
    port map (
            O => \N__22531\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__22528\,
            I => \N__22525\
        );

    \I__2981\ : InMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__2979\ : Span4Mux_v
    port map (
            O => \N__22519\,
            I => \N__22515\
        );

    \I__2978\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22512\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__22515\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__22512\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__2975\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22504\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__22498\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__2971\ : InMux
    port map (
            O => \N__22495\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__2970\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22489\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__22489\,
            I => \N__22486\
        );

    \I__2968\ : Span4Mux_v
    port map (
            O => \N__22486\,
            I => \N__22482\
        );

    \I__2967\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22479\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__22482\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__22479\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__2964\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22471\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22468\
        );

    \I__2962\ : Span4Mux_h
    port map (
            O => \N__22468\,
            I => \N__22465\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__22465\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__2960\ : InMux
    port map (
            O => \N__22462\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__2959\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__22453\,
            I => \N__22449\
        );

    \I__2956\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22446\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__22449\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__22446\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__2953\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22438\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22435\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__22432\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__2949\ : InMux
    port map (
            O => \N__22429\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__22420\,
            I => \N__22416\
        );

    \I__2945\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22413\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__22416\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__22413\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__22405\,
            I => \N__22402\
        );

    \I__2940\ : Span4Mux_h
    port map (
            O => \N__22402\,
            I => \N__22399\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__22399\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22396\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22393\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22390\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__2935\ : InMux
    port map (
            O => \N__22387\,
            I => \bfn_7_14_0_\
        );

    \I__2934\ : InMux
    port map (
            O => \N__22384\,
            I => \N__22381\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__22381\,
            I => \N__22378\
        );

    \I__2932\ : Odrv12
    port map (
            O => \N__22378\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_0\
        );

    \I__2931\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22372\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__22372\,
            I => \N__22369\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__22369\,
            I => \N__22366\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__22366\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_5\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__22363\,
            I => \N__22360\
        );

    \I__2926\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__2924\ : Span4Mux_h
    port map (
            O => \N__22354\,
            I => \N__22351\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__22351\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__2921\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__2919\ : Span4Mux_v
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__22336\,
            I => \N__22333\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__22333\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__2915\ : InMux
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__22324\,
            I => \N__22321\
        );

    \I__2913\ : Span4Mux_h
    port map (
            O => \N__22321\,
            I => \N__22318\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__22318\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__22315\,
            I => \N__22312\
        );

    \I__2910\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22309\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22309\,
            I => \N__22306\
        );

    \I__2908\ : Span4Mux_h
    port map (
            O => \N__22306\,
            I => \N__22303\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__22303\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__22300\,
            I => \N__22297\
        );

    \I__2905\ : InMux
    port map (
            O => \N__22297\,
            I => \N__22293\
        );

    \I__2904\ : InMux
    port map (
            O => \N__22296\,
            I => \N__22290\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22287\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__22290\,
            I => \N__22283\
        );

    \I__2901\ : Span4Mux_v
    port map (
            O => \N__22287\,
            I => \N__22280\
        );

    \I__2900\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22277\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__22283\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__22280\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__22277\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__22270\,
            I => \N__22267\
        );

    \I__2895\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22264\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__22264\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__22261\,
            I => \N__22258\
        );

    \I__2892\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22255\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__22255\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__22252\,
            I => \N__22249\
        );

    \I__2889\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22246\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__22246\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__22243\,
            I => \N__22240\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__22237\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__22234\,
            I => \N__22231\
        );

    \I__2883\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__22228\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__22225\,
            I => \N__22222\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22219\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22219\,
            I => \N__22216\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__22216\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__22213\,
            I => \N__22210\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22210\,
            I => \N__22207\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__22207\,
            I => \N__22204\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__22204\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__22201\,
            I => \N__22194\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__22200\,
            I => \N__22190\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__22199\,
            I => \N__22186\
        );

    \I__2870\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22171\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22197\,
            I => \N__22171\
        );

    \I__2868\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22171\
        );

    \I__2867\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22171\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22171\
        );

    \I__2865\ : InMux
    port map (
            O => \N__22189\,
            I => \N__22171\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22171\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22168\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__22168\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__22165\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22159\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__22159\,
            I => \current_shift_inst.PI_CTRL.un1_enablelt3_0\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__22156\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__22153\,
            I => \N__22150\
        );

    \I__2856\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22147\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__22147\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22141\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__22132\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22126\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__22126\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__22123\,
            I => \N__22120\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22117\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__22117\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__22114\,
            I => \N__22111\
        );

    \I__2843\ : InMux
    port map (
            O => \N__22111\,
            I => \N__22108\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__22108\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22102\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__22102\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22096\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__22096\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22093\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22087\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22087\,
            I => \N__22084\
        );

    \I__2834\ : Odrv12
    port map (
            O => \N__22084\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__22081\,
            I => \N__22078\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22078\,
            I => \N__22075\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__22075\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__22072\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22066\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__22066\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__2827\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22060\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22054\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__22054\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__2823\ : InMux
    port map (
            O => \N__22051\,
            I => \N__22048\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22048\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22045\,
            I => \N__22042\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__22042\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22036\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22036\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__22033\,
            I => \N__22030\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22030\,
            I => \N__22027\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__22027\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__22021\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22015\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22015\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__22012\,
            I => \N__22009\
        );

    \I__2809\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__22003\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21997\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__21997\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__21994\,
            I => \N__21991\
        );

    \I__2803\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21988\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21985\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__21985\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__2800\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21979\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__21979\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__21976\,
            I => \N__21973\
        );

    \I__2797\ : InMux
    port map (
            O => \N__21973\,
            I => \N__21970\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__21970\,
            I => \N__21967\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__21967\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__2794\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21961\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__21961\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__21958\,
            I => \N__21955\
        );

    \I__2791\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21952\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__21952\,
            I => \N__21949\
        );

    \I__2789\ : Odrv12
    port map (
            O => \N__21949\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__2788\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21943\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__21943\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__21940\,
            I => \N__21937\
        );

    \I__2785\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21934\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__21934\,
            I => \N__21931\
        );

    \I__2783\ : Span4Mux_h
    port map (
            O => \N__21931\,
            I => \N__21928\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__21928\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__2781\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21922\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__21922\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__2779\ : InMux
    port map (
            O => \N__21919\,
            I => \N__21916\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__21916\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__2777\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21910\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__21910\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__21907\,
            I => \N__21904\
        );

    \I__2774\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21901\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__21901\,
            I => \N__21898\
        );

    \I__2772\ : Span4Mux_h
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__21895\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__2770\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__21889\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__2768\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__21880\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__21877\,
            I => \un2_counter_5_cascade_\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__21874\,
            I => \N__21869\
        );

    \I__2763\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21866\
        );

    \I__2762\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21860\
        );

    \I__2761\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21860\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21857\
        );

    \I__2759\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21854\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__21860\,
            I => \counterZ0Z_0\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__21857\,
            I => \counterZ0Z_0\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__21854\,
            I => \counterZ0Z_0\
        );

    \I__2755\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21843\
        );

    \I__2754\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21840\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__21843\,
            I => \counterZ0Z_11\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__21840\,
            I => \counterZ0Z_11\
        );

    \I__2751\ : InMux
    port map (
            O => \N__21835\,
            I => \N__21831\
        );

    \I__2750\ : InMux
    port map (
            O => \N__21834\,
            I => \N__21828\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__21831\,
            I => \counterZ0Z_9\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__21828\,
            I => \counterZ0Z_9\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__21823\,
            I => \N__21819\
        );

    \I__2746\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21816\
        );

    \I__2745\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21813\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__21816\,
            I => \counterZ0Z_12\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__21813\,
            I => \counterZ0Z_12\
        );

    \I__2742\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21804\
        );

    \I__2741\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21801\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21798\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__21801\,
            I => \counterZ0Z_8\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__21798\,
            I => \counterZ0Z_8\
        );

    \I__2737\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21787\
        );

    \I__2736\ : InMux
    port map (
            O => \N__21792\,
            I => \N__21782\
        );

    \I__2735\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21779\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21776\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21773\
        );

    \I__2732\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21770\
        );

    \I__2731\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21767\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__21782\,
            I => \N__21760\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__21779\,
            I => \N__21760\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__21776\,
            I => \N__21760\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__21773\,
            I => un2_counter_7
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__21770\,
            I => un2_counter_7
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__21767\,
            I => un2_counter_7
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__21760\,
            I => un2_counter_7
        );

    \I__2723\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21741\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21741\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21736\
        );

    \I__2720\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21736\
        );

    \I__2719\ : InMux
    port map (
            O => \N__21747\,
            I => \N__21733\
        );

    \I__2718\ : InMux
    port map (
            O => \N__21746\,
            I => \N__21730\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__21741\,
            I => un2_counter_8
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__21736\,
            I => un2_counter_8
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__21733\,
            I => un2_counter_8
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__21730\,
            I => un2_counter_8
        );

    \I__2713\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21711\
        );

    \I__2712\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21711\
        );

    \I__2711\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21706\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21706\
        );

    \I__2709\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21703\
        );

    \I__2708\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21700\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__21711\,
            I => un2_counter_9
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__21706\,
            I => un2_counter_9
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__21703\,
            I => un2_counter_9
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__21700\,
            I => un2_counter_9
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__21691\,
            I => \N__21686\
        );

    \I__2702\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21683\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__21689\,
            I => \N__21679\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21676\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21673\
        );

    \I__2698\ : InMux
    port map (
            O => \N__21682\,
            I => \N__21670\
        );

    \I__2697\ : InMux
    port map (
            O => \N__21679\,
            I => \N__21667\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__21676\,
            I => clk_10khz_i
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__21673\,
            I => clk_10khz_i
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__21670\,
            I => clk_10khz_i
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21667\,
            I => clk_10khz_i
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__21658\,
            I => \N__21654\
        );

    \I__2691\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21651\
        );

    \I__2690\ : InMux
    port map (
            O => \N__21654\,
            I => \N__21648\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__21651\,
            I => \counterZ0Z_6\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__21648\,
            I => \counterZ0Z_6\
        );

    \I__2687\ : InMux
    port map (
            O => \N__21643\,
            I => un5_counter_cry_5
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__2685\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21634\,
            I => \counter_RNO_0Z0Z_7\
        );

    \I__2683\ : InMux
    port map (
            O => \N__21631\,
            I => un5_counter_cry_6
        );

    \I__2682\ : InMux
    port map (
            O => \N__21628\,
            I => un5_counter_cry_7
        );

    \I__2681\ : InMux
    port map (
            O => \N__21625\,
            I => \bfn_5_8_0_\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__21622\,
            I => \N__21619\
        );

    \I__2679\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__21616\,
            I => \counter_RNO_0Z0Z_10\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21613\,
            I => un5_counter_cry_9
        );

    \I__2676\ : InMux
    port map (
            O => \N__21610\,
            I => un5_counter_cry_10
        );

    \I__2675\ : InMux
    port map (
            O => \N__21607\,
            I => un5_counter_cry_11
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__21604\,
            I => \N__21601\
        );

    \I__2673\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21598\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__21598\,
            I => \counter_RNO_0Z0Z_12\
        );

    \I__2671\ : InMux
    port map (
            O => \N__21595\,
            I => \N__21591\
        );

    \I__2670\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21588\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__21591\,
            I => \counterZ0Z_10\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__21588\,
            I => \counterZ0Z_10\
        );

    \I__2667\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21579\
        );

    \I__2666\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21576\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__21579\,
            I => \counterZ0Z_7\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__21576\,
            I => \counterZ0Z_7\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21567\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21564\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__21567\,
            I => \N__21561\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21564\,
            I => \counterZ0Z_2\
        );

    \I__2659\ : Odrv12
    port map (
            O => \N__21561\,
            I => \counterZ0Z_2\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__21556\,
            I => \N__21553\
        );

    \I__2657\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21549\
        );

    \I__2656\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21545\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21542\
        );

    \I__2654\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21539\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__21545\,
            I => \counterZ0Z_1\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__21542\,
            I => \counterZ0Z_1\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__21539\,
            I => \counterZ0Z_1\
        );

    \I__2650\ : InMux
    port map (
            O => \N__21532\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__21529\,
            I => \N__21523\
        );

    \I__2648\ : InMux
    port map (
            O => \N__21528\,
            I => \N__21518\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__21527\,
            I => \N__21515\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \N__21509\
        );

    \I__2645\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21506\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21500\
        );

    \I__2643\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21500\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21497\
        );

    \I__2641\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21494\
        );

    \I__2640\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21485\
        );

    \I__2639\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21485\
        );

    \I__2638\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21485\
        );

    \I__2637\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21485\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21482\
        );

    \I__2635\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21479\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__21500\,
            I => \N__21476\
        );

    \I__2633\ : Span12Mux_s7_v
    port map (
            O => \N__21497\,
            I => \N__21469\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__21494\,
            I => \N__21469\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__21485\,
            I => \N__21469\
        );

    \I__2630\ : Span4Mux_h
    port map (
            O => \N__21482\,
            I => \N__21466\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21463\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__21476\,
            I => \N__21460\
        );

    \I__2627\ : Span12Mux_v
    port map (
            O => \N__21469\,
            I => \N__21457\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__21466\,
            I => \N__21454\
        );

    \I__2625\ : Span12Mux_s4_h
    port map (
            O => \N__21463\,
            I => \N__21451\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__21460\,
            I => \N__21448\
        );

    \I__2623\ : Odrv12
    port map (
            O => \N__21457\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__21454\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__21451\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__21448\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21436\
        );

    \I__2618\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21433\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__21433\,
            I => \N__21430\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__21430\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__21427\,
            I => \N__21424\
        );

    \I__2614\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21421\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21418\
        );

    \I__2612\ : Odrv4
    port map (
            O => \N__21418\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2611\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21412\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__21412\,
            I => \N__21409\
        );

    \I__2609\ : Span4Mux_s2_v
    port map (
            O => \N__21409\,
            I => \N__21406\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__21406\,
            I => un7_start_stop_0_a3
        );

    \I__2607\ : InMux
    port map (
            O => \N__21403\,
            I => un5_counter_cry_1
        );

    \I__2606\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21396\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21399\,
            I => \N__21393\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__21396\,
            I => \counterZ0Z_3\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__21393\,
            I => \counterZ0Z_3\
        );

    \I__2602\ : InMux
    port map (
            O => \N__21388\,
            I => un5_counter_cry_2
        );

    \I__2601\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21381\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21378\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__21381\,
            I => \counterZ0Z_4\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__21378\,
            I => \counterZ0Z_4\
        );

    \I__2597\ : InMux
    port map (
            O => \N__21373\,
            I => un5_counter_cry_3
        );

    \I__2596\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21366\
        );

    \I__2595\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21363\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__21366\,
            I => \counterZ0Z_5\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__21363\,
            I => \counterZ0Z_5\
        );

    \I__2592\ : InMux
    port map (
            O => \N__21358\,
            I => un5_counter_cry_4
        );

    \I__2591\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21351\
        );

    \I__2590\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21348\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21345\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__21348\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__21345\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2586\ : InMux
    port map (
            O => \N__21340\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2585\ : InMux
    port map (
            O => \N__21337\,
            I => \N__21333\
        );

    \I__2584\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21330\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__21333\,
            I => \N__21325\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__21330\,
            I => \N__21325\
        );

    \I__2581\ : Span4Mux_h
    port map (
            O => \N__21325\,
            I => \N__21322\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__21322\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21319\,
            I => \bfn_4_20_0_\
        );

    \I__2578\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21312\
        );

    \I__2577\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21309\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21312\,
            I => \N__21306\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__21309\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__21306\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21301\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\
        );

    \I__2572\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21292\
        );

    \I__2571\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21292\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__21292\,
            I => \N__21289\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__21289\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2568\ : InMux
    port map (
            O => \N__21286\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2567\ : InMux
    port map (
            O => \N__21283\,
            I => \N__21280\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21280\,
            I => \N__21276\
        );

    \I__2565\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21273\
        );

    \I__2564\ : Odrv4
    port map (
            O => \N__21276\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__21273\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21268\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2561\ : InMux
    port map (
            O => \N__21265\,
            I => \N__21262\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__21262\,
            I => \N__21258\
        );

    \I__2559\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21255\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__21258\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__21255\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21250\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2555\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21243\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21240\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__21243\,
            I => \N__21235\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21240\,
            I => \N__21235\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__21235\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2550\ : InMux
    port map (
            O => \N__21232\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__2548\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21222\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21219\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21216\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21219\,
            I => \N__21211\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__21216\,
            I => \N__21211\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__21211\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2542\ : InMux
    port map (
            O => \N__21208\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21205\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21196\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21193\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__21193\,
            I => \N__21190\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__21190\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__21187\,
            I => \N__21184\
        );

    \I__2534\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21180\
        );

    \I__2533\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21177\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__21180\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__21177\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2530\ : InMux
    port map (
            O => \N__21172\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2529\ : InMux
    port map (
            O => \N__21169\,
            I => \N__21166\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__21166\,
            I => \N__21163\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__21163\,
            I => \N__21159\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21156\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__21159\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21156\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2523\ : InMux
    port map (
            O => \N__21151\,
            I => \bfn_4_19_0_\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__21148\,
            I => \N__21145\
        );

    \I__2521\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21142\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N__21139\
        );

    \I__2519\ : Odrv4
    port map (
            O => \N__21139\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__21136\,
            I => \N__21133\
        );

    \I__2517\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21130\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21126\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21123\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__21126\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21123\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21118\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21111\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__21114\,
            I => \N__21108\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21111\,
            I => \N__21105\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21102\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__21105\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21102\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2505\ : InMux
    port map (
            O => \N__21097\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21088\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21088\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__21088\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21085\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__21082\,
            I => \N__21079\
        );

    \I__2499\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21073\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21078\,
            I => \N__21073\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__21073\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21070\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21063\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21060\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21063\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21060\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21055\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__21052\,
            I => \N__21048\
        );

    \I__2489\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21043\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21048\,
            I => \N__21043\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21043\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2486\ : InMux
    port map (
            O => \N__21040\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__21037\,
            I => \N__21034\
        );

    \I__2484\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21030\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21026\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__21030\,
            I => \N__21023\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21029\,
            I => \N__21020\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21017\
        );

    \I__2479\ : Span4Mux_h
    port map (
            O => \N__21023\,
            I => \N__21012\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__21020\,
            I => \N__21012\
        );

    \I__2477\ : Span4Mux_h
    port map (
            O => \N__21017\,
            I => \N__21009\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__21012\,
            I => \N__21006\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__21009\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__21006\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21001\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__20998\,
            I => \N__20995\
        );

    \I__2471\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20991\
        );

    \I__2470\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20987\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__20991\,
            I => \N__20984\
        );

    \I__2468\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20981\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20978\
        );

    \I__2466\ : Span4Mux_h
    port map (
            O => \N__20984\,
            I => \N__20973\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20973\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__20978\,
            I => \N__20970\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__20973\,
            I => \N__20967\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__20970\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__20967\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2460\ : InMux
    port map (
            O => \N__20962\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__20959\,
            I => \N__20956\
        );

    \I__2458\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20953\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20949\
        );

    \I__2456\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20946\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__20949\,
            I => \N__20942\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20939\
        );

    \I__2453\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20936\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__20942\,
            I => \N__20933\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__20939\,
            I => \N__20930\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20927\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__20933\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__20930\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2447\ : Odrv12
    port map (
            O => \N__20927\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2446\ : InMux
    port map (
            O => \N__20920\,
            I => \bfn_4_18_0_\
        );

    \I__2445\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20914\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20911\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__20911\,
            I => \N__20907\
        );

    \I__2442\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20904\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__20907\,
            I => \N__20900\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__20904\,
            I => \N__20897\
        );

    \I__2439\ : InMux
    port map (
            O => \N__20903\,
            I => \N__20894\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__20900\,
            I => \N__20891\
        );

    \I__2437\ : Span4Mux_h
    port map (
            O => \N__20897\,
            I => \N__20888\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20885\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__20891\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__20888\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2433\ : Odrv12
    port map (
            O => \N__20885\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2432\ : InMux
    port map (
            O => \N__20878\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__20875\,
            I => \N__20871\
        );

    \I__2430\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20868\
        );

    \I__2429\ : InMux
    port map (
            O => \N__20871\,
            I => \N__20865\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__20868\,
            I => \N__20860\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20860\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__20860\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2425\ : InMux
    port map (
            O => \N__20857\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2424\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20851\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__20851\,
            I => \N__20847\
        );

    \I__2422\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20844\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__20847\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__20844\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2419\ : InMux
    port map (
            O => \N__20839\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2418\ : InMux
    port map (
            O => \N__20836\,
            I => \N__20830\
        );

    \I__2417\ : InMux
    port map (
            O => \N__20835\,
            I => \N__20830\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__20830\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2415\ : InMux
    port map (
            O => \N__20827\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2414\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20817\
        );

    \I__2412\ : InMux
    port map (
            O => \N__20820\,
            I => \N__20814\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__20817\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__20814\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2409\ : InMux
    port map (
            O => \N__20809\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2408\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20800\
        );

    \I__2407\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20800\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__20800\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__20797\,
            I => \N__20794\
        );

    \I__2404\ : InMux
    port map (
            O => \N__20794\,
            I => \N__20791\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__20791\,
            I => \N__20788\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__20788\,
            I => \N__20785\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__20785\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__20782\,
            I => \N__20779\
        );

    \I__2399\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20776\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__2397\ : Span4Mux_h
    port map (
            O => \N__20773\,
            I => \N__20770\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__20770\,
            I => \N__20767\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__20767\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__20764\,
            I => \N__20761\
        );

    \I__2393\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20758\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20755\
        );

    \I__2391\ : Span4Mux_h
    port map (
            O => \N__20755\,
            I => \N__20752\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__2389\ : Odrv4
    port map (
            O => \N__20749\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2388\ : InMux
    port map (
            O => \N__20746\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__20743\,
            I => \N__20740\
        );

    \I__2386\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20737\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__20737\,
            I => \N__20734\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__20734\,
            I => \N__20731\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__20731\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__20728\,
            I => \N__20725\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20722\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__2379\ : Span4Mux_v
    port map (
            O => \N__20719\,
            I => \N__20716\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__20713\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2376\ : InMux
    port map (
            O => \N__20710\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2375\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20703\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__20706\,
            I => \N__20700\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__20703\,
            I => \N__20696\
        );

    \I__2372\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20693\
        );

    \I__2371\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20690\
        );

    \I__2370\ : Span4Mux_h
    port map (
            O => \N__20696\,
            I => \N__20687\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20682\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__20690\,
            I => \N__20682\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__20687\,
            I => \N__20677\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__20682\,
            I => \N__20677\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__20677\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2364\ : InMux
    port map (
            O => \N__20674\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__20671\,
            I => \N__20668\
        );

    \I__2362\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20664\
        );

    \I__2361\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20661\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20656\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__20661\,
            I => \N__20653\
        );

    \I__2358\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20650\
        );

    \I__2357\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20647\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__20656\,
            I => \N__20638\
        );

    \I__2355\ : Span4Mux_s2_h
    port map (
            O => \N__20653\,
            I => \N__20638\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20638\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20647\,
            I => \N__20638\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__20638\,
            I => \N__20635\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__20635\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20632\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2349\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20625\
        );

    \I__2348\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20621\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__20625\,
            I => \N__20618\
        );

    \I__2346\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20615\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__20621\,
            I => \N__20612\
        );

    \I__2344\ : Span12Mux_s4_h
    port map (
            O => \N__20618\,
            I => \N__20607\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__20615\,
            I => \N__20607\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__20612\,
            I => \N__20604\
        );

    \I__2341\ : Odrv12
    port map (
            O => \N__20607\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__20604\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2339\ : InMux
    port map (
            O => \N__20599\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__20596\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__20593\,
            I => \N__20590\
        );

    \I__2336\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20586\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20583\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20580\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__20583\,
            I => \N__20577\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__20580\,
            I => \N__20574\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__20577\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__20574\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2329\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20566\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20562\
        );

    \I__2327\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20559\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__20562\,
            I => \clk_10khz_RNIIENAZ0Z2\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__20559\,
            I => \clk_10khz_RNIIENAZ0Z2\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20551\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20551\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\
        );

    \I__2322\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20545\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__20545\,
            I => \N__20542\
        );

    \I__2320\ : Glb2LocalMux
    port map (
            O => \N__20542\,
            I => \N__20539\
        );

    \I__2319\ : GlobalMux
    port map (
            O => \N__20539\,
            I => clk_12mhz
        );

    \I__2318\ : IoInMux
    port map (
            O => \N__20536\,
            I => \N__20533\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__20533\,
            I => \N__20530\
        );

    \I__2316\ : Span4Mux_s0_v
    port map (
            O => \N__20530\,
            I => \N__20527\
        );

    \I__2315\ : Span4Mux_h
    port map (
            O => \N__20527\,
            I => \N__20524\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__20524\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2313\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20518\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__20518\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_8\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__20515\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20509\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__20509\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__20506\,
            I => \N__20503\
        );

    \I__2307\ : InMux
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__20500\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__20497\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__2304\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20491\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__20491\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__2302\ : InMux
    port map (
            O => \N__20488\,
            I => \N__20485\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__20485\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__2300\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__20476\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__20473\,
            I => \N__20470\
        );

    \I__2296\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20464\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__20464\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__2293\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__20458\,
            I => \N__20455\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__20455\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__2290\ : InMux
    port map (
            O => \N__20452\,
            I => \N__20449\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__20449\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\
        );

    \I__2288\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__20443\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__20437\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\
        );

    \I__2284\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20431\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__20431\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\
        );

    \I__2282\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__20425\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\
        );

    \I__2280\ : InMux
    port map (
            O => \N__20422\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19\
        );

    \I__2279\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20416\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__20416\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20410\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20410\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20404\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__20404\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2273\ : InMux
    port map (
            O => \N__20401\,
            I => \N__20398\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__20398\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__2270\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20388\
        );

    \I__2269\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20385\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__20388\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__20385\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20380\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_6\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__20374\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__20371\,
            I => \N__20368\
        );

    \I__2262\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20365\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__20365\,
            I => \N__20362\
        );

    \I__2260\ : Span4Mux_s3_h
    port map (
            O => \N__20362\,
            I => \N__20359\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__20359\,
            I => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\
        );

    \I__2258\ : InMux
    port map (
            O => \N__20356\,
            I => \bfn_3_13_0_\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20350\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20350\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\
        );

    \I__2255\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20344\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__20344\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\
        );

    \I__2253\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20338\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__20338\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20332\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__20332\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20329\,
            I => \N__20326\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__20326\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\
        );

    \I__2247\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20320\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__20320\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\
        );

    \I__2245\ : InMux
    port map (
            O => \N__20317\,
            I => \N__20312\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \N__20309\
        );

    \I__2243\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20306\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20303\
        );

    \I__2241\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20300\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__20306\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__20303\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__20300\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_12\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20293\,
            I => \N__20289\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20292\,
            I => \N__20286\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20283\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__20286\,
            I => \N__20280\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__20283\,
            I => \N__20275\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__20280\,
            I => \N__20275\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__20275\,
            I => \pwm_generator_inst.un3_threshold_acc\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20269\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20266\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__20263\,
            I => \pwm_generator_inst.O_12\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20257\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__20257\,
            I => \N__20253\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20250\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__20253\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__20250\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\
        );

    \I__2221\ : InMux
    port map (
            O => \N__20245\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_0\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__2219\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20236\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__20236\,
            I => \N__20233\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__20233\,
            I => \N__20230\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__20230\,
            I => \pwm_generator_inst.O_13\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20220\
        );

    \I__2213\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20217\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__20220\,
            I => \N__20212\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__20217\,
            I => \N__20212\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__20212\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\
        );

    \I__2209\ : InMux
    port map (
            O => \N__20209\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_1\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20203\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__20203\,
            I => \N__20200\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__20197\,
            I => \pwm_generator_inst.O_14\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__20194\,
            I => \N__20191\
        );

    \I__2203\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20187\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20184\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__20187\,
            I => \N__20179\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__20184\,
            I => \N__20179\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__20179\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20176\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_2\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20173\,
            I => \N__20170\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__20170\,
            I => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__20167\,
            I => \N__20164\
        );

    \I__2194\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20161\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20157\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20154\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__20157\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__20154\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20149\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_3\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__20146\,
            I => \N__20143\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20140\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__20140\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20131\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20131\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__20131\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20128\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_4\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20122\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20122\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\
        );

    \I__2179\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20115\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20112\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__20115\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__20112\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20107\,
            I => \pwm_generator_inst.un3_threshold_acc_cry_5\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20099\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20096\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20093\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__20099\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__20096\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__20093\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_14\
        );

    \I__2168\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20083\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20083\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20080\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_13\
        );

    \I__2165\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20074\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__20074\,
            I => \N__20071\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__20071\,
            I => \N__20068\
        );

    \I__2162\ : Odrv4
    port map (
            O => \N__20068\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20065\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_14\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20058\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20055\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__20058\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20055\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20047\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__20047\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20044\,
            I => \bfn_3_11_0_\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__20041\,
            I => \N__20038\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20035\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20035\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20032\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_16\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20026\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20023\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_17\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20020\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18\
        );

    \I__2145\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__20014\,
            I => \N__20011\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__20011\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\
        );

    \I__2142\ : InMux
    port map (
            O => \N__20008\,
            I => \N__20004\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20000\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__19997\
        );

    \I__2139\ : InMux
    port map (
            O => \N__20003\,
            I => \N__19994\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20000\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__19997\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__19994\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_15\
        );

    \I__2135\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19982\
        );

    \I__2134\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19977\
        );

    \I__2133\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19977\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19974\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__19977\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__19974\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_18\
        );

    \I__2129\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19964\
        );

    \I__2128\ : InMux
    port map (
            O => \N__19968\,
            I => \N__19959\
        );

    \I__2127\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19959\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__19964\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__19959\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_17\
        );

    \I__2124\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__19948\,
            I => \N__19945\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__19945\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2120\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__19939\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_7\
        );

    \I__2118\ : InMux
    port map (
            O => \N__19936\,
            I => \N__19933\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__19930\,
            I => \N__19927\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__19927\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2114\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19921\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__19921\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_8\
        );

    \I__2112\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19915\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19912\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__19909\,
            I => \pwm_generator_inst.O_9\
        );

    \I__2108\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__19903\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_9\
        );

    \I__2106\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19897\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19892\
        );

    \I__2104\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19889\
        );

    \I__2103\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19886\
        );

    \I__2102\ : Span4Mux_h
    port map (
            O => \N__19892\,
            I => \N__19883\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__19889\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__19886\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__19883\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_10\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__19876\,
            I => \N__19873\
        );

    \I__2097\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19870\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__19867\,
            I => \N__19864\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__19864\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\
        );

    \I__2093\ : InMux
    port map (
            O => \N__19861\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_9\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__19858\,
            I => \N__19854\
        );

    \I__2091\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19842\
        );

    \I__2090\ : InMux
    port map (
            O => \N__19854\,
            I => \N__19839\
        );

    \I__2089\ : InMux
    port map (
            O => \N__19853\,
            I => \N__19828\
        );

    \I__2088\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19828\
        );

    \I__2087\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19828\
        );

    \I__2086\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19828\
        );

    \I__2085\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19828\
        );

    \I__2084\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19825\
        );

    \I__2083\ : InMux
    port map (
            O => \N__19847\,
            I => \N__19818\
        );

    \I__2082\ : InMux
    port map (
            O => \N__19846\,
            I => \N__19818\
        );

    \I__2081\ : InMux
    port map (
            O => \N__19845\,
            I => \N__19818\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__19842\,
            I => \N__19811\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__19839\,
            I => \N__19811\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__19828\,
            I => \N__19811\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19807\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__19818\,
            I => \N__19802\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__19811\,
            I => \N__19802\
        );

    \I__2074\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19799\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__19807\,
            I => \N__19796\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__19802\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__19799\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__19796\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\
        );

    \I__2069\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19786\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19783\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__19783\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_1\
        );

    \I__2066\ : InMux
    port map (
            O => \N__19780\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_10\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__19777\,
            I => \N__19774\
        );

    \I__2064\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__19771\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\
        );

    \I__2062\ : InMux
    port map (
            O => \N__19768\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_11\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__19765\,
            I => \N__19760\
        );

    \I__2060\ : InMux
    port map (
            O => \N__19764\,
            I => \N__19757\
        );

    \I__2059\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19754\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19751\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__19757\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__19754\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__19751\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_13\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__19741\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\
        );

    \I__2052\ : InMux
    port map (
            O => \N__19738\,
            I => \pwm_generator_inst.un15_threshold_acc_1_cry_12\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19722\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19722\
        );

    \I__2049\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19717\
        );

    \I__2048\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19717\
        );

    \I__2047\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19706\
        );

    \I__2046\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19706\
        );

    \I__2045\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19706\
        );

    \I__2044\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19706\
        );

    \I__2043\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19706\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__19722\,
            I => \N__19699\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19699\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19696\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19693\
        );

    \I__2038\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19690\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__19699\,
            I => \N__19687\
        );

    \I__2036\ : Span4Mux_h
    port map (
            O => \N__19696\,
            I => \N__19684\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19693\,
            I => \N__19681\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__19690\,
            I => pwm_duty_input_6
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__19687\,
            I => pwm_duty_input_6
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__19684\,
            I => pwm_duty_input_6
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__19681\,
            I => pwm_duty_input_6
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__19672\,
            I => \N__19666\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__19671\,
            I => \N__19663\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__19670\,
            I => \N__19660\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19649\
        );

    \I__2026\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19649\
        );

    \I__2025\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19644\
        );

    \I__2024\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19644\
        );

    \I__2023\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19641\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19658\,
            I => \N__19630\
        );

    \I__2021\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19630\
        );

    \I__2020\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19630\
        );

    \I__2019\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19630\
        );

    \I__2018\ : InMux
    port map (
            O => \N__19654\,
            I => \N__19630\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19649\,
            I => \N__19627\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__19644\,
            I => \N__19624\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__19641\,
            I => i8_mux
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__19630\,
            I => i8_mux
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__19627\,
            I => i8_mux
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__19624\,
            I => i8_mux
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__19615\,
            I => \N__19604\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__19614\,
            I => \N__19601\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__19613\,
            I => \N__19598\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__19612\,
            I => \N__19595\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__19611\,
            I => \N__19592\
        );

    \I__2006\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19587\
        );

    \I__2005\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19587\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19582\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19582\
        );

    \I__2002\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19574\
        );

    \I__2001\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19574\
        );

    \I__2000\ : InMux
    port map (
            O => \N__19598\,
            I => \N__19574\
        );

    \I__1999\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19569\
        );

    \I__1998\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19569\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__19587\,
            I => \N__19564\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__19582\,
            I => \N__19564\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19561\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__19574\,
            I => \N__19556\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__19569\,
            I => \N__19556\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__19564\,
            I => \N__19553\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__19561\,
            I => \N__19548\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__19556\,
            I => \N__19548\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__19553\,
            I => \N__19545\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__19548\,
            I => \N_28_mux\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__19545\,
            I => \N_28_mux\
        );

    \I__1986\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19537\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__19537\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\
        );

    \I__1984\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19531\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__19531\,
            I => \N__19528\
        );

    \I__1982\ : Span4Mux_v
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__19525\,
            I => \pwm_generator_inst.O_0\
        );

    \I__1980\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19519\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__19519\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_0\
        );

    \I__1978\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19513\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19510\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__19510\,
            I => \N__19507\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__19507\,
            I => \pwm_generator_inst.O_1\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19501\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_1\
        );

    \I__1972\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19495\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__19495\,
            I => \N__19492\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__19492\,
            I => \N__19489\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__19489\,
            I => \pwm_generator_inst.O_2\
        );

    \I__1968\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__19483\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_2\
        );

    \I__1966\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19477\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__19474\,
            I => \N__19471\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__19471\,
            I => \pwm_generator_inst.O_3\
        );

    \I__1962\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19465\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__19465\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_3\
        );

    \I__1960\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19459\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__19456\,
            I => \N__19453\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__19453\,
            I => \pwm_generator_inst.O_4\
        );

    \I__1956\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19447\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__19447\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_4\
        );

    \I__1954\ : InMux
    port map (
            O => \N__19444\,
            I => \N__19441\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__19438\,
            I => \N__19435\
        );

    \I__1951\ : Odrv4
    port map (
            O => \N__19435\,
            I => \pwm_generator_inst.O_5\
        );

    \I__1950\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19429\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__19429\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_5\
        );

    \I__1948\ : InMux
    port map (
            O => \N__19426\,
            I => \N__19423\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__1946\ : Span4Mux_h
    port map (
            O => \N__19420\,
            I => \N__19417\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__19417\,
            I => \pwm_generator_inst.O_6\
        );

    \I__1944\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__19411\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_6\
        );

    \I__1942\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__19405\,
            I => \N__19402\
        );

    \I__1940\ : Span4Mux_s2_v
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__19399\,
            I => \N_22_i_i\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__19393\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__1935\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19384\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__19384\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\
        );

    \I__1933\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19378\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__19378\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_6\
        );

    \I__1931\ : InMux
    port map (
            O => \N__19375\,
            I => \N__19372\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__19372\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\
        );

    \I__1929\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__19366\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\
        );

    \I__1927\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19360\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__19360\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\
        );

    \I__1925\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__19354\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\
        );

    \I__1923\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19348\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__19348\,
            I => \N__19344\
        );

    \I__1921\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19341\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__19344\,
            I => \N__19336\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__19341\,
            I => \N__19336\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__19336\,
            I => \pwm_generator_inst.O_10\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19330\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19327\
        );

    \I__1915\ : Odrv12
    port map (
            O => \N__19327\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_0\
        );

    \I__1914\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19321\,
            I => \N__19318\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__19318\,
            I => \N__19314\
        );

    \I__1911\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19311\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__19314\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__19311\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__19306\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1907\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19300\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__19300\,
            I => \N__19295\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19292\
        );

    \I__1904\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19289\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__19295\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__19292\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__19289\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__1900\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19278\
        );

    \I__1899\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19271\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19268\
        );

    \I__1897\ : InMux
    port map (
            O => \N__19277\,
            I => \N__19259\
        );

    \I__1896\ : InMux
    port map (
            O => \N__19276\,
            I => \N__19259\
        );

    \I__1895\ : InMux
    port map (
            O => \N__19275\,
            I => \N__19259\
        );

    \I__1894\ : InMux
    port map (
            O => \N__19274\,
            I => \N__19259\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__19271\,
            I => \N__19251\
        );

    \I__1892\ : Span4Mux_s2_h
    port map (
            O => \N__19268\,
            I => \N__19251\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19259\,
            I => \N__19251\
        );

    \I__1890\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19248\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__19251\,
            I => \N__19243\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__19248\,
            I => \N__19243\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__19243\,
            I => \current_shift_inst.PI_CTRL.N_118\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__19240\,
            I => \N__19236\
        );

    \I__1885\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19229\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19218\
        );

    \I__1883\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19218\
        );

    \I__1882\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19218\
        );

    \I__1881\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19218\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19218\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19229\,
            I => \N__19213\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__19218\,
            I => \N__19210\
        );

    \I__1877\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19207\
        );

    \I__1876\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19204\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__19213\,
            I => \N__19194\
        );

    \I__1874\ : Span4Mux_s2_h
    port map (
            O => \N__19210\,
            I => \N__19194\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19194\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__19204\,
            I => \N__19194\
        );

    \I__1871\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19191\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__19194\,
            I => \N__19186\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__19191\,
            I => \N__19186\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__19186\,
            I => \current_shift_inst.PI_CTRL.N_178\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__19183\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19177\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19177\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__1864\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19171\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__19171\,
            I => \N__19168\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__19168\,
            I => \N__19165\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__19165\,
            I => \N__19162\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__19162\,
            I => \pwm_generator_inst.un2_threshold_acc_2_11\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19159\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__19156\,
            I => \N__19153\
        );

    \I__1857\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19150\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__19150\,
            I => \N__19147\
        );

    \I__1855\ : Span4Mux_h
    port map (
            O => \N__19147\,
            I => \N__19144\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__19141\,
            I => \pwm_generator_inst.un2_threshold_acc_2_12\
        );

    \I__1852\ : InMux
    port map (
            O => \N__19138\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19132\,
            I => \N__19129\
        );

    \I__1849\ : Span4Mux_h
    port map (
            O => \N__19129\,
            I => \N__19126\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__19126\,
            I => \N__19123\
        );

    \I__1847\ : Odrv4
    port map (
            O => \N__19123\,
            I => \pwm_generator_inst.un2_threshold_acc_2_13\
        );

    \I__1846\ : InMux
    port map (
            O => \N__19120\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__19117\,
            I => \N__19114\
        );

    \I__1844\ : InMux
    port map (
            O => \N__19114\,
            I => \N__19111\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__1842\ : Span4Mux_h
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__19102\,
            I => \pwm_generator_inst.un2_threshold_acc_2_14\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19099\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\
        );

    \I__1838\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__19087\,
            I => \N__19084\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__19084\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\
        );

    \I__1833\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__19078\,
            I => \N__19071\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19068\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__19076\,
            I => \N__19065\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__19075\,
            I => \N__19061\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__19074\,
            I => \N__19057\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__19071\,
            I => \N__19051\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__19068\,
            I => \N__19051\
        );

    \I__1825\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19038\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19038\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19061\,
            I => \N__19038\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19038\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19038\
        );

    \I__1820\ : InMux
    port map (
            O => \N__19056\,
            I => \N__19038\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__19051\,
            I => \N__19035\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__19038\,
            I => \N__19032\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__19035\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__19032\,
            I => \pwm_generator_inst.un2_threshold_acc_1_25\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19027\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\
        );

    \I__1814\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19021\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__19021\,
            I => \N__19018\
        );

    \I__1812\ : Span4Mux_v
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__19015\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19012\,
            I => \bfn_2_14_0_\
        );

    \I__1809\ : InMux
    port map (
            O => \N__19009\,
            I => \N__19006\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__19006\,
            I => \N__19001\
        );

    \I__1807\ : InMux
    port map (
            O => \N__19005\,
            I => \N__18996\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19004\,
            I => \N__18996\
        );

    \I__1805\ : Span4Mux_s2_h
    port map (
            O => \N__19001\,
            I => \N__18991\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__18996\,
            I => \N__18991\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__18991\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1802\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18985\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__18985\,
            I => \current_shift_inst.PI_CTRL.N_98\
        );

    \I__1800\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__1799\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18976\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18971\
        );

    \I__1797\ : InMux
    port map (
            O => \N__18975\,
            I => \N__18966\
        );

    \I__1796\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18966\
        );

    \I__1795\ : Span4Mux_s2_h
    port map (
            O => \N__18971\,
            I => \N__18960\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__18966\,
            I => \N__18960\
        );

    \I__1793\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18957\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__18960\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__18957\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1790\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18949\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__18949\,
            I => \N__18946\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__18946\,
            I => \pwm_generator_inst.un2_threshold_acc_1_18\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__18943\,
            I => \N__18940\
        );

    \I__1786\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18937\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__18937\,
            I => \N__18934\
        );

    \I__1784\ : Span4Mux_h
    port map (
            O => \N__18934\,
            I => \N__18931\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__18931\,
            I => \N__18928\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__18928\,
            I => \pwm_generator_inst.un2_threshold_acc_2_3\
        );

    \I__1781\ : InMux
    port map (
            O => \N__18925\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\
        );

    \I__1780\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18919\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__18919\,
            I => \N__18916\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__18916\,
            I => \pwm_generator_inst.un2_threshold_acc_1_19\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__18913\,
            I => \N__18910\
        );

    \I__1776\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18907\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18904\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__18904\,
            I => \N__18901\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__18901\,
            I => \N__18898\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__18898\,
            I => \pwm_generator_inst.un2_threshold_acc_2_4\
        );

    \I__1771\ : InMux
    port map (
            O => \N__18895\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\
        );

    \I__1770\ : InMux
    port map (
            O => \N__18892\,
            I => \N__18889\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__18889\,
            I => \N__18886\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__18886\,
            I => \N__18883\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__18883\,
            I => \N__18880\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__18880\,
            I => \pwm_generator_inst.un2_threshold_acc_2_5\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__18877\,
            I => \N__18874\
        );

    \I__1764\ : InMux
    port map (
            O => \N__18874\,
            I => \N__18871\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__18871\,
            I => \N__18868\
        );

    \I__1762\ : Odrv4
    port map (
            O => \N__18868\,
            I => \pwm_generator_inst.un2_threshold_acc_1_20\
        );

    \I__1761\ : InMux
    port map (
            O => \N__18865\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\
        );

    \I__1760\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18859\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__18859\,
            I => \N__18856\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__18856\,
            I => \N__18853\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__18853\,
            I => \N__18850\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__18850\,
            I => \pwm_generator_inst.un2_threshold_acc_2_6\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__18847\,
            I => \N__18844\
        );

    \I__1754\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18841\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18838\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__18838\,
            I => \pwm_generator_inst.un2_threshold_acc_1_21\
        );

    \I__1751\ : InMux
    port map (
            O => \N__18835\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\
        );

    \I__1750\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18829\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__18829\,
            I => \N__18826\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__18826\,
            I => \N__18823\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__18823\,
            I => \N__18820\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__18820\,
            I => \pwm_generator_inst.un2_threshold_acc_2_7\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__18817\,
            I => \N__18814\
        );

    \I__1744\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18811\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__18811\,
            I => \N__18808\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__18808\,
            I => \pwm_generator_inst.un2_threshold_acc_1_22\
        );

    \I__1741\ : InMux
    port map (
            O => \N__18805\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\
        );

    \I__1740\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18799\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__18799\,
            I => \N__18796\
        );

    \I__1738\ : Span4Mux_h
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__18793\,
            I => \pwm_generator_inst.un2_threshold_acc_1_23\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__18790\,
            I => \N__18787\
        );

    \I__1735\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18784\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__18784\,
            I => \N__18781\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__18781\,
            I => \N__18778\
        );

    \I__1732\ : Span4Mux_v
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__18775\,
            I => \pwm_generator_inst.un2_threshold_acc_2_8\
        );

    \I__1730\ : InMux
    port map (
            O => \N__18772\,
            I => \bfn_2_13_0_\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18766\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__18766\,
            I => \N__18763\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__18763\,
            I => \pwm_generator_inst.un2_threshold_acc_1_24\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__18760\,
            I => \N__18757\
        );

    \I__1725\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18754\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__18754\,
            I => \N__18751\
        );

    \I__1723\ : Span4Mux_v
    port map (
            O => \N__18751\,
            I => \N__18748\
        );

    \I__1722\ : Span4Mux_v
    port map (
            O => \N__18748\,
            I => \N__18745\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__18745\,
            I => \pwm_generator_inst.un2_threshold_acc_2_9\
        );

    \I__1720\ : InMux
    port map (
            O => \N__18742\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__18739\,
            I => \N__18736\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18733\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18730\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__18730\,
            I => \N__18727\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__18727\,
            I => \N__18724\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__18724\,
            I => \pwm_generator_inst.un2_threshold_acc_2_10\
        );

    \I__1713\ : InMux
    port map (
            O => \N__18721\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__18718\,
            I => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\
        );

    \I__1711\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18712\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__18712\,
            I => \N__18709\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__18709\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_6\
        );

    \I__1708\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__18703\,
            I => \N__18700\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__18700\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_7\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__18697\,
            I => \N__18694\
        );

    \I__1704\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18691\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__18691\,
            I => \N__18688\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__18688\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_8\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__18679\,
            I => \N__18676\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__18676\,
            I => \N__18673\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__18673\,
            I => \pwm_generator_inst.un2_threshold_acc_2_0\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__18670\,
            I => \N__18667\
        );

    \I__1695\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18664\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__18664\,
            I => \N__18661\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__18661\,
            I => \N__18658\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__18658\,
            I => \pwm_generator_inst.un2_threshold_acc_1_15\
        );

    \I__1691\ : InMux
    port map (
            O => \N__18655\,
            I => \N__18652\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__18652\,
            I => \N__18649\
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__18649\,
            I => \pwm_generator_inst.un2_threshold_acc_1_16\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__18646\,
            I => \N__18643\
        );

    \I__1687\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18640\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__18637\,
            I => \N__18634\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__18634\,
            I => \N__18631\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__18631\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1\
        );

    \I__1682\ : InMux
    port map (
            O => \N__18628\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18622\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__18622\,
            I => \N__18619\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__18619\,
            I => \pwm_generator_inst.un2_threshold_acc_1_17\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__18616\,
            I => \N__18613\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18610\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__18607\,
            I => \N__18604\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__18601\,
            I => \pwm_generator_inst.un2_threshold_acc_2_2\
        );

    \I__1672\ : InMux
    port map (
            O => \N__18598\,
            I => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\
        );

    \I__1671\ : InMux
    port map (
            O => \N__18595\,
            I => \bfn_2_9_0_\
        );

    \I__1670\ : InMux
    port map (
            O => \N__18592\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_8\
        );

    \I__1669\ : InMux
    port map (
            O => \N__18589\,
            I => \N__18586\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__18586\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_4\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__18583\,
            I => \N__18579\
        );

    \I__1666\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18576\
        );

    \I__1665\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18572\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__18576\,
            I => \N__18569\
        );

    \I__1663\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18566\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__18572\,
            I => \N__18563\
        );

    \I__1661\ : Span4Mux_s1_h
    port map (
            O => \N__18569\,
            I => \N__18560\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__18566\,
            I => pwm_duty_input_8
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__18563\,
            I => pwm_duty_input_8
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__18560\,
            I => pwm_duty_input_8
        );

    \I__1657\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18524\
        );

    \I__1656\ : InMux
    port map (
            O => \N__18552\,
            I => \N__18524\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18551\,
            I => \N__18524\
        );

    \I__1654\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18524\
        );

    \I__1653\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18524\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18524\
        );

    \I__1651\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18524\
        );

    \I__1650\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18524\
        );

    \I__1649\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18519\
        );

    \I__1648\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18519\
        );

    \I__1647\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18513\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__18542\,
            I => \N__18510\
        );

    \I__1645\ : InMux
    port map (
            O => \N__18541\,
            I => \N__18507\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__18524\,
            I => \N__18504\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__18519\,
            I => \N__18501\
        );

    \I__1642\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18494\
        );

    \I__1641\ : InMux
    port map (
            O => \N__18517\,
            I => \N__18494\
        );

    \I__1640\ : InMux
    port map (
            O => \N__18516\,
            I => \N__18494\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__18513\,
            I => \N__18491\
        );

    \I__1638\ : InMux
    port map (
            O => \N__18510\,
            I => \N__18488\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__18507\,
            I => \N__18471\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__18504\,
            I => \N__18471\
        );

    \I__1635\ : Span4Mux_s1_h
    port map (
            O => \N__18501\,
            I => \N__18471\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__18494\,
            I => \N__18471\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__18491\,
            I => \N__18466\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__18488\,
            I => \N__18466\
        );

    \I__1631\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18463\
        );

    \I__1630\ : InMux
    port map (
            O => \N__18486\,
            I => \N__18448\
        );

    \I__1629\ : InMux
    port map (
            O => \N__18485\,
            I => \N__18448\
        );

    \I__1628\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18448\
        );

    \I__1627\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18448\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18448\
        );

    \I__1625\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18448\
        );

    \I__1624\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18448\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__18471\,
            I => \N__18445\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__18466\,
            I => pwm_duty_input_10
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__18463\,
            I => pwm_duty_input_10
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__18448\,
            I => pwm_duty_input_10
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__18445\,
            I => pwm_duty_input_10
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__18436\,
            I => \N__18433\
        );

    \I__1617\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18427\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__18427\,
            I => \current_shift_inst.PI_CTRL.m7_2\
        );

    \I__1614\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18419\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18416\
        );

    \I__1612\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18413\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18410\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__18416\,
            I => \N__18407\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__18413\,
            I => pwm_duty_input_7
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__18410\,
            I => pwm_duty_input_7
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__18407\,
            I => pwm_duty_input_7
        );

    \I__1606\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18397\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__18397\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_5\
        );

    \I__1604\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18391\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__18391\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_2\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__18388\,
            I => \N__18385\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18382\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__18382\,
            I => \pwm_generator_inst.un19_threshold_acc_axb_3\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__18379\,
            I => \N__18376\
        );

    \I__1598\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18373\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__18373\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\
        );

    \I__1596\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18367\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__18367\,
            I => \pwm_generator_inst.threshold_ACCZ0Z_9\
        );

    \I__1594\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18361\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__18361\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\
        );

    \I__1592\ : InMux
    port map (
            O => \N__18358\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__18355\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_1\
        );

    \I__1590\ : InMux
    port map (
            O => \N__18352\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_2\
        );

    \I__1589\ : InMux
    port map (
            O => \N__18349\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_3\
        );

    \I__1588\ : InMux
    port map (
            O => \N__18346\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_4\
        );

    \I__1587\ : InMux
    port map (
            O => \N__18343\,
            I => \N__18340\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__18340\,
            I => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\
        );

    \I__1585\ : InMux
    port map (
            O => \N__18337\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_5\
        );

    \I__1584\ : InMux
    port map (
            O => \N__18334\,
            I => \pwm_generator_inst.un19_threshold_acc_cry_6\
        );

    \I__1583\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18327\
        );

    \I__1582\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18324\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__18327\,
            I => pwm_duty_input_2
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__18324\,
            I => pwm_duty_input_2
        );

    \I__1579\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18314\
        );

    \I__1578\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18311\
        );

    \I__1577\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18308\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__18314\,
            I => \N__18305\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18302\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18297\
        );

    \I__1573\ : Span4Mux_s1_h
    port map (
            O => \N__18305\,
            I => \N__18297\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__18302\,
            I => pwm_duty_input_3
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__18297\,
            I => pwm_duty_input_3
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__18292\,
            I => \N__18289\
        );

    \I__1569\ : InMux
    port map (
            O => \N__18289\,
            I => \N__18285\
        );

    \I__1568\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18282\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__18285\,
            I => pwm_duty_input_0
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__18282\,
            I => pwm_duty_input_0
        );

    \I__1565\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18273\
        );

    \I__1564\ : InMux
    port map (
            O => \N__18276\,
            I => \N__18270\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__18273\,
            I => \N__18267\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__18270\,
            I => \N__18264\
        );

    \I__1561\ : Span4Mux_v
    port map (
            O => \N__18267\,
            I => \N__18261\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__18264\,
            I => pwm_duty_input_1
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__18261\,
            I => pwm_duty_input_1
        );

    \I__1558\ : InMux
    port map (
            O => \N__18256\,
            I => \N__18253\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__18253\,
            I => \N__18250\
        );

    \I__1556\ : Odrv12
    port map (
            O => \N__18250\,
            I => \current_shift_inst.PI_CTRL.m14_2\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__18247\,
            I => \current_shift_inst.PI_CTRL.N_19_cascade_\
        );

    \I__1554\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18240\
        );

    \I__1553\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18236\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18233\
        );

    \I__1551\ : InMux
    port map (
            O => \N__18239\,
            I => \N__18230\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__18236\,
            I => pwm_duty_input_4
        );

    \I__1549\ : Odrv12
    port map (
            O => \N__18233\,
            I => pwm_duty_input_4
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18230\,
            I => pwm_duty_input_4
        );

    \I__1547\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18220\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__18217\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__1544\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18209\
        );

    \I__1543\ : InMux
    port map (
            O => \N__18213\,
            I => \N__18204\
        );

    \I__1542\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18204\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__18209\,
            I => \N__18199\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__18204\,
            I => \N__18199\
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__18199\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1538\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18193\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__18193\,
            I => \N__18189\
        );

    \I__1536\ : InMux
    port map (
            O => \N__18192\,
            I => \N__18186\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__18189\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__18186\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_15\
        );

    \I__1533\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18178\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__18178\,
            I => \pwm_generator_inst.un2_threshold_acc_2_1_16\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__18175\,
            I => \N__18171\
        );

    \I__1530\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18167\
        );

    \I__1529\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18162\
        );

    \I__1528\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18162\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__18167\,
            I => \N__18159\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__18162\,
            I => pwm_duty_input_9
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__18159\,
            I => pwm_duty_input_9
        );

    \I__1524\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18147\
        );

    \I__1523\ : InMux
    port map (
            O => \N__18153\,
            I => \N__18147\
        );

    \I__1522\ : InMux
    port map (
            O => \N__18152\,
            I => \N__18144\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__18147\,
            I => \N__18141\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18138\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__18141\,
            I => pwm_duty_input_5
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__18138\,
            I => pwm_duty_input_5
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_6\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_14\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_10_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_22\,
            carryinitout => \bfn_10_24_0_\
        );

    \IN_MUX_bfv_10_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_0_cry_30\,
            carryinitout => \bfn_10_25_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_counter_cry_8,
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            carryinitout => \bfn_3_14_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_18_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_8_0_\
        );

    \IN_MUX_bfv_18_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_18_9_0_\
        );

    \IN_MUX_bfv_18_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_18_10_0_\
        );

    \IN_MUX_bfv_12_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_24_0_\
        );

    \IN_MUX_bfv_12_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_12_25_0_\
        );

    \IN_MUX_bfv_12_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_12_26_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_8\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_16\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_5_cry_24\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_3_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_9_0_\
        );

    \IN_MUX_bfv_3_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            carryinitout => \bfn_3_10_0_\
        );

    \IN_MUX_bfv_3_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            carryinitout => \bfn_3_11_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_10_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_12_0_\
        );

    \IN_MUX_bfv_10_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_10_13_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_13_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_21_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_18_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_23_0_\
        );

    \IN_MUX_bfv_18_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_18_24_0_\
        );

    \IN_MUX_bfv_18_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_18_25_0_\
        );

    \IN_MUX_bfv_18_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_18_26_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_17_25_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_7\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_15\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_14_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.z_cry_23\,
            carryinitout => \bfn_14_21_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_8\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_16\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_cry_24\,
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_16_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_17_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_17_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_17_14_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_16_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_23_0_\
        );

    \IN_MUX_bfv_16_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_24_0_\
        );

    \IN_MUX_bfv_16_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_25_0_\
        );

    \IN_MUX_bfv_14_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_22_0_\
        );

    \IN_MUX_bfv_14_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_7\,
            carryinitout => \bfn_14_23_0_\
        );

    \IN_MUX_bfv_14_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_15\,
            carryinitout => \bfn_14_24_0_\
        );

    \IN_MUX_bfv_14_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_phase.counter_cry_23\,
            carryinitout => \bfn_14_25_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_11_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_7\,
            carryinitout => \bfn_11_21_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_15\,
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_1_cry_23\,
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_4_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryinitout => \bfn_4_19_0_\
        );

    \IN_MUX_bfv_4_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryinitout => \bfn_4_20_0_\
        );

    \IN_MUX_bfv_8_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_17_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryinitout => \bfn_8_19_0_\
        );

    \IN_MUX_bfv_8_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryinitout => \bfn_8_20_0_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27256\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_336_i_g\
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__23056\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_187_i_g\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__30070\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_phase.N_188_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__43350\,
            CLKHFEN => \N__43449\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__43493\,
            RGB2PWM => \N__19408\,
            RGB1 => rgb_g_wire,
            CURREN => \N__43334\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__21415\,
            RGB0PWM => \N__48279\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__19081\,
            in1 => \N__18192\,
            in2 => \_gnd_net_\,
            in3 => \N__18487\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21528\,
            lcout => pwm_duty_input_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48874\,
            ce => \N__25133\,
            sr => \N__48174\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIDE9T_3_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__18318\,
            in1 => \N__18244\,
            in2 => \N__18175\,
            in3 => \N__18154\,
            lcout => \current_shift_inst.PI_CTRL.m7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNILM9T_5_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18170\,
            in1 => \N__18424\,
            in2 => \N__18583\,
            in3 => \N__18153\,
            lcout => \current_shift_inst.PI_CTRL.m14_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__18196\,
            in1 => \N__19077\,
            in2 => \N__18542\,
            in3 => \N__18181\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001110"
        )
    port map (
            in0 => \N__20917\,
            in1 => \N__19239\,
            in2 => \N__21527\,
            in3 => \N__19282\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48871\,
            ce => \N__25081\,
            sr => \N__48202\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19235\,
            in1 => \N__21514\,
            in2 => \N__20959\,
            in3 => \N__19277\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48868\,
            ce => \N__25132\,
            sr => \N__48209\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001100"
        )
    port map (
            in0 => \N__19274\,
            in1 => \N__20629\,
            in2 => \N__21526\,
            in3 => \N__19232\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48868\,
            ce => \N__25132\,
            sr => \N__48209\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19234\,
            in1 => \N__21513\,
            in2 => \N__20998\,
            in3 => \N__19276\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48868\,
            ce => \N__25132\,
            sr => \N__48209\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011011101"
        )
    port map (
            in0 => \N__18982\,
            in1 => \N__20707\,
            in2 => \N__19240\,
            in3 => \N__19324\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48868\,
            ce => \N__25132\,
            sr => \N__48209\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19233\,
            in1 => \N__21512\,
            in2 => \N__21037\,
            in3 => \N__19275\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48868\,
            ce => \N__25132\,
            sr => \N__48209\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18214\,
            in1 => \N__18981\,
            in2 => \N__20764\,
            in3 => \N__19009\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48868\,
            ce => \N__25132\,
            sr => \N__48209\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18975\,
            in1 => \N__18213\,
            in2 => \N__20728\,
            in3 => \N__19005\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48864\,
            ce => \N__25077\,
            sr => \N__48213\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__18974\,
            in1 => \N__18212\,
            in2 => \N__20782\,
            in3 => \N__19004\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48864\,
            ce => \N__25077\,
            sr => \N__48213\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__20589\,
            in1 => \N__18223\,
            in2 => \N__20671\,
            in3 => \N__19281\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48864\,
            ce => \N__25077\,
            sr => \N__48213\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIUU8T_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__18331\,
            in1 => \N__18317\,
            in2 => \N__18292\,
            in3 => \N__18276\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIK2D32_4_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__18256\,
            in1 => \N__18541\,
            in2 => \N__18247\,
            in3 => \N__18243\,
            lcout => \N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19896\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19347\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__20667\,
            in1 => \N__19303\,
            in2 => \N__21529\,
            in3 => \N__19216\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20659\,
            in2 => \_gnd_net_\,
            in3 => \N__20699\,
            lcout => \current_shift_inst.PI_CTRL.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21505\,
            in1 => \N__19299\,
            in2 => \_gnd_net_\,
            in3 => \N__19203\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_6_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__19610\,
            in1 => \N__19734\,
            in2 => \N__19671\,
            in3 => \N__18343\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48873\,
            ce => 'H',
            sr => \N__48175\
        );

    \pwm_generator_inst.threshold_ACC_1_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__19609\,
            in1 => \N__18364\,
            in2 => \N__19670\,
            in3 => \N__19735\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48873\,
            ce => 'H',
            sr => \N__48175\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19333\,
            in2 => \N__19858\,
            in3 => \N__19857\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19789\,
            in2 => \_gnd_net_\,
            in3 => \N__18358\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18394\,
            in2 => \_gnd_net_\,
            in3 => \N__18355\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18388\,
            in3 => \N__18352\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18589\,
            in2 => \_gnd_net_\,
            in3 => \N__18349\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18400\,
            in2 => \_gnd_net_\,
            in3 => \N__18346\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18715\,
            in2 => \_gnd_net_\,
            in3 => \N__18337\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18706\,
            in2 => \_gnd_net_\,
            in3 => \N__18334\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18697\,
            in3 => \N__18595\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => \pwm_generator_inst.un19_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__20017\,
            in1 => \N__19853\,
            in2 => \N__20371\,
            in3 => \N__18592\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__19851\,
            in1 => \N__20086\,
            in2 => \N__20194\,
            in3 => \N__20103\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNIVCED1_7_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__18575\,
            in1 => \N__18543\,
            in2 => \N__18436\,
            in3 => \N__18422\,
            lcout => i8_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__19852\,
            in1 => \N__20077\,
            in2 => \N__20167\,
            in3 => \N__20008\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20260\,
            in1 => \N__20317\,
            in2 => \N__19777\,
            in3 => \N__19850\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__19849\,
            in1 => \N__19744\,
            in2 => \N__20227\,
            in3 => \N__19763\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_9_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000000110000"
        )
    port map (
            in0 => \N__19581\,
            in1 => \N__19659\,
            in2 => \N__18379\,
            in3 => \N__19704\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48865\,
            ce => 'H',
            sr => \N__48203\
        );

    \pwm_generator_inst.threshold_9_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18370\,
            lcout => \pwm_generator_inst.thresholdZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48865\,
            ce => 'H',
            sr => \N__48203\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20223\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20190\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20136\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_16\,
            ltout => \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20137\,
            in1 => \N__20050\,
            in2 => \N__18718\,
            in3 => \N__19845\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__20119\,
            in1 => \N__19969\,
            in2 => \N__20041\,
            in3 => \N__19846\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__19987\,
            in1 => \N__19847\,
            in2 => \N__20395\,
            in3 => \N__20029\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_axb_4_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18685\,
            in2 => \N__18670\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18655\,
            in2 => \N__18646\,
            in3 => \N__18628\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18625\,
            in2 => \N__18616\,
            in3 => \N__18598\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18952\,
            in2 => \N__18943\,
            in3 => \N__18925\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18922\,
            in2 => \N__18913\,
            in3 => \N__18895\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18892\,
            in2 => \N__18877\,
            in3 => \N__18865\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18862\,
            in2 => \N__18847\,
            in3 => \N__18835\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18832\,
            in2 => \N__18817\,
            in3 => \N__18805\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18802\,
            in2 => \N__18790\,
            in3 => \N__18772\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18769\,
            in2 => \N__18760\,
            in3 => \N__18742\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19056\,
            in2 => \N__18739\,
            in3 => \N__18721\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19174\,
            in2 => \N__19074\,
            in3 => \N__19159\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19060\,
            in2 => \N__19156\,
            in3 => \N__19138\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19135\,
            in2 => \N__19075\,
            in3 => \N__19120\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19064\,
            in2 => \N__19117\,
            in3 => \N__19099\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19096\,
            in2 => \N__19076\,
            in3 => \N__19027\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_acc_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_acc_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__20419\,
            in1 => \N__19024\,
            in2 => \_gnd_net_\,
            in3 => \N__19012\,
            lcout => \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__19317\,
            in1 => \N__19217\,
            in2 => \N__20706\,
            in3 => \N__18965\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__18988\,
            in1 => \N__21522\,
            in2 => \N__20593\,
            in3 => \N__19258\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__19895\,
            in1 => \N__19351\,
            in2 => \N__19876\,
            in3 => \N__19810\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__20660\,
            in1 => \N__21521\,
            in2 => \_gnd_net_\,
            in3 => \N__19298\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20628\,
            in2 => \_gnd_net_\,
            in3 => \N__20994\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20952\,
            in1 => \N__21033\,
            in2 => \N__19306\,
            in3 => \N__20910\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20461\,
            in1 => \N__20512\,
            in2 => \N__20506\,
            in3 => \N__20488\,
            lcout => \current_shift_inst.PI_CTRL.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_10_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20407\,
            in1 => \N__20482\,
            in2 => \N__20473\,
            in3 => \N__19180\,
            lcout => \current_shift_inst.PI_CTRL.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20824\,
            in2 => \_gnd_net_\,
            in3 => \N__21169\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISHP8_10_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20413\,
            in1 => \N__20854\,
            in2 => \N__19183\,
            in3 => \N__20874\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28105\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48801\,
            ce => \N__25152\,
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28762\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48801\,
            ce => \N__25152\,
            sr => \N__48238\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28684\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48801\,
            ce => \N__25152\,
            sr => \N__48238\
        );

    \current_shift_inst.N_22_i_i_LC_2_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__48278\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31032\,
            lcout => \N_22_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_7_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__19732\,
            in1 => \N__19608\,
            in2 => \N__19672\,
            in3 => \N__19396\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48872\,
            ce => 'H',
            sr => \N__48163\
        );

    \pwm_generator_inst.threshold_ACC_0_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__19607\,
            in1 => \N__19733\,
            in2 => \N__19390\,
            in3 => \N__19669\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48872\,
            ce => 'H',
            sr => \N__48163\
        );

    \pwm_generator_inst.threshold_6_LC_3_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19381\,
            lcout => \pwm_generator_inst.thresholdZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48872\,
            ce => 'H',
            sr => \N__48163\
        );

    \pwm_generator_inst.threshold_ACC_4_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__19728\,
            in1 => \N__19657\,
            in2 => \N__19614\,
            in3 => \N__19375\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48869\,
            ce => 'H',
            sr => \N__48176\
        );

    \pwm_generator_inst.threshold_ACC_2_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__19654\,
            in1 => \N__19730\,
            in2 => \N__19611\,
            in3 => \N__19369\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48869\,
            ce => 'H',
            sr => \N__48176\
        );

    \pwm_generator_inst.threshold_ACC_3_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__19727\,
            in1 => \N__19656\,
            in2 => \N__19613\,
            in3 => \N__19363\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48869\,
            ce => 'H',
            sr => \N__48176\
        );

    \pwm_generator_inst.threshold_ACC_8_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__19655\,
            in1 => \N__19731\,
            in2 => \N__19612\,
            in3 => \N__19357\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48869\,
            ce => 'H',
            sr => \N__48176\
        );

    \pwm_generator_inst.threshold_ACC_5_LC_3_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__19729\,
            in1 => \N__19658\,
            in2 => \N__19615\,
            in3 => \N__19540\,
            lcout => \pwm_generator_inst.threshold_ACCZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48869\,
            ce => 'H',
            sr => \N__48176\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19522\,
            in2 => \_gnd_net_\,
            in3 => \N__19534\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_3_9_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19504\,
            in2 => \_gnd_net_\,
            in3 => \N__19516\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19486\,
            in2 => \_gnd_net_\,
            in3 => \N__19498\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19468\,
            in2 => \_gnd_net_\,
            in3 => \N__19480\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19450\,
            in2 => \_gnd_net_\,
            in3 => \N__19462\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19432\,
            in2 => \_gnd_net_\,
            in3 => \N__19444\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19414\,
            in2 => \_gnd_net_\,
            in3 => \N__19426\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19942\,
            in2 => \_gnd_net_\,
            in3 => \N__19954\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19924\,
            in2 => \_gnd_net_\,
            in3 => \N__19936\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_3_10_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19906\,
            in2 => \_gnd_net_\,
            in3 => \N__19918\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19900\,
            in2 => \_gnd_net_\,
            in3 => \N__19861\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__19848\,
            in1 => \N__20293\,
            in2 => \_gnd_net_\,
            in3 => \N__19780\,
            lcout => \pwm_generator_inst.un19_threshold_acc_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20316\,
            in3 => \N__19768\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19765\,
            in3 => \N__19738\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20102\,
            in2 => \_gnd_net_\,
            in3 => \N__20080\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20003\,
            in2 => \_gnd_net_\,
            in3 => \N__20065\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20061\,
            in2 => \_gnd_net_\,
            in3 => \N__20044\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_3_11_0_\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19967\,
            in2 => \_gnd_net_\,
            in3 => \N__20032\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19985\,
            in2 => \_gnd_net_\,
            in3 => \N__20023\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_acc_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_acc_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20020\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20160\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19986\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20391\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__19968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20118\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__20315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20256\,
            lcout => \pwm_generator_inst.un15_threshold_acc_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20292\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20272\,
            in2 => \_gnd_net_\,
            in3 => \N__20245\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20242\,
            in3 => \N__20209\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20206\,
            in2 => \_gnd_net_\,
            in3 => \N__20176\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20173\,
            in2 => \_gnd_net_\,
            in3 => \N__20149\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43430\,
            in2 => \N__20146\,
            in3 => \N__20128\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20125\,
            in2 => \N__43472\,
            in3 => \N__20107\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20401\,
            in2 => \N__43434\,
            in3 => \N__20380\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20377\,
            in2 => \_gnd_net_\,
            in3 => \N__20356\,
            lcout => \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20353\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20347\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20341\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20335\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20329\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20323\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20452\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20446\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_14_0_\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20440\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20434\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20428\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_acc_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_acc_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20422\,
            lcout => \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIEE4_12_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21247\,
            in1 => \N__20806\,
            in2 => \N__21229\,
            in3 => \N__20836\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_0_10_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26376\,
            in1 => \N__26338\,
            in2 => \N__26301\,
            in3 => \N__26257\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_8_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRMD4_17_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21337\,
            in1 => \N__21115\,
            in2 => \N__21136\,
            in3 => \N__21298\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMJ62_12_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20835\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIU8H5_14_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20805\,
            in1 => \N__21297\,
            in2 => \N__20515\,
            in3 => \N__21336\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_10_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21246\,
            in1 => \N__20850\,
            in2 => \N__20875\,
            in3 => \N__21225\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21129\,
            in1 => \N__21162\,
            in2 => \N__21114\,
            in3 => \N__21183\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPM62_13_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21316\,
            in2 => \_gnd_net_\,
            in3 => \N__20820\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIKAQ8_27_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21265\,
            in1 => \N__21283\,
            in2 => \N__20497\,
            in3 => \N__20494\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI9LI5_19_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21094\,
            in1 => \N__20554\,
            in2 => \N__21082\,
            in3 => \N__21315\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIEAE4_15_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21067\,
            in1 => \N__21354\,
            in2 => \N__21187\,
            in3 => \N__21051\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21066\,
            in1 => \N__21078\,
            in2 => \N__21052\,
            in3 => \N__21093\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1082_27_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21261\,
            in2 => \_gnd_net_\,
            in3 => \N__21279\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20548\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNII76D_3_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21369\,
            in1 => \N__21384\,
            in2 => \N__21658\,
            in3 => \N__21399\,
            lcout => un2_counter_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_7_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__21721\,
            in1 => \N__21751\,
            in2 => \N__21640\,
            in3 => \N__21786\,
            lcout => \counterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48866\,
            ce => 'H',
            sr => \N__48164\
        );

    \counter_12_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__21750\,
            in1 => \N__21785\,
            in2 => \N__21604\,
            in3 => \N__21720\,
            lcout => \counterZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48866\,
            ce => 'H',
            sr => \N__48164\
        );

    \counter_1_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21552\,
            in2 => \_gnd_net_\,
            in3 => \N__21872\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48860\,
            ce => 'H',
            sr => \N__48177\
        );

    \pwm_generator_inst.threshold_8_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20521\,
            lcout => \pwm_generator_inst.thresholdZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48860\,
            ce => 'H',
            sr => \N__48177\
        );

    \counter_10_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__21719\,
            in1 => \N__21749\,
            in2 => \N__21622\,
            in3 => \N__21792\,
            lcout => \counterZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48860\,
            ce => 'H',
            sr => \N__48177\
        );

    \counter_0_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__21748\,
            in1 => \N__21791\,
            in2 => \N__21874\,
            in3 => \N__21718\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48860\,
            ce => 'H',
            sr => \N__48177\
        );

    \clk_10khz_RNIIENA2_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__21746\,
            in1 => \N__21790\,
            in2 => \N__21689\,
            in3 => \N__21716\,
            lcout => \clk_10khz_RNIIENAZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__30988\,
            in1 => \N__21682\,
            in2 => \_gnd_net_\,
            in3 => \N__20565\,
            lcout => \N_717_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIU1LD_7_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20903\,
            in2 => \_gnd_net_\,
            in3 => \N__20990\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20945\,
            in1 => \N__21029\,
            in2 => \N__20596\,
            in3 => \N__20624\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.phase_valid_RNISLOR2_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21690\,
            in1 => \N__24277\,
            in2 => \N__31033\,
            in3 => \N__20569\,
            lcout => \current_shift_inst.phase_valid_RNISLORZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23368\,
            in1 => \N__23492\,
            in2 => \N__23632\,
            in3 => \N__22507\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23365\,
            in1 => \N__23483\,
            in2 => \N__23629\,
            in3 => \N__22753\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010001010"
        )
    port map (
            in0 => \N__22726\,
            in1 => \N__23493\,
            in2 => \N__23391\,
            in3 => \N__23613\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23366\,
            in1 => \N__23484\,
            in2 => \N__23630\,
            in3 => \N__22699\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__23369\,
            in1 => \N__23617\,
            in2 => \N__23502\,
            in3 => \N__22669\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23367\,
            in1 => \N__23488\,
            in2 => \N__23631\,
            in3 => \N__22642\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__23370\,
            in1 => \N__23621\,
            in2 => \N__23503\,
            in3 => \N__22612\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48829\,
            ce => 'H',
            sr => \N__48214\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28183\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48819\,
            ce => \N__25054\,
            sr => \N__48218\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23938\,
            in2 => \N__20797\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23914\,
            in2 => \N__22138\,
            in3 => \N__20746\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23889\,
            in2 => \N__20743\,
            in3 => \N__20710\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23845\,
            in2 => \N__22123\,
            in3 => \N__20674\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22144\,
            in2 => \N__23818\,
            in3 => \N__20632\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23769\,
            in2 => \N__22081\,
            in3 => \N__20599\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23731\,
            in2 => \N__23002\,
            in3 => \N__21001\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23695\,
            in2 => \N__22153\,
            in3 => \N__20962\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__48802\,
            ce => \N__25106\,
            sr => \N__48225\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24079\,
            in2 => \N__22969\,
            in3 => \N__20920\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24034\,
            in2 => \N__22114\,
            in3 => \N__20878\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26256\,
            in2 => \N__22252\,
            in3 => \N__20857\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26574\,
            in2 => \N__22225\,
            in3 => \N__20839\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26784\,
            in2 => \N__22939\,
            in3 => \N__20827\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26653\,
            in2 => \N__21439\,
            in3 => \N__20809\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_4_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22129\,
            in2 => \N__26695\,
            in3 => \N__21205\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26337\,
            in2 => \N__21202\,
            in3 => \N__21172\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__48792\,
            ce => \N__25154\,
            sr => \N__48230\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26612\,
            in2 => \N__22270\,
            in3 => \N__21151\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_4_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24826\,
            in2 => \N__21148\,
            in3 => \N__21118\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24184\,
            in2 => \N__21427\,
            in3 => \N__21097\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24937\,
            in2 => \N__22261\,
            in3 => \N__21085\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24972\,
            in2 => \N__22984\,
            in3 => \N__21070\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26407\,
            in2 => \N__22243\,
            in3 => \N__21055\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24883\,
            in2 => \N__22234\,
            in3 => \N__21040\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26375\,
            in2 => \N__22213\,
            in3 => \N__21340\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__48784\,
            ce => \N__25064\,
            sr => \N__48233\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26490\,
            in2 => \N__22954\,
            in3 => \N__21319\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_4_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_4_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26530\,
            in2 => \N__22199\,
            in3 => \N__21301\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22189\,
            in2 => \N__26455\,
            in3 => \N__21286\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26819\,
            in2 => \N__22200\,
            in3 => \N__21268\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_4_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22193\,
            in2 => \N__26749\,
            in3 => \N__21250\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26294\,
            in2 => \N__22201\,
            in3 => \N__21232\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22197\,
            in2 => \N__26191\,
            in3 => \N__21208\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22198\,
            in1 => \N__25520\,
            in2 => \_gnd_net_\,
            in3 => \N__21532\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48775\,
            ce => \N__25155\,
            sr => \N__48236\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_4_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28212\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48766\,
            ce => \N__25172\,
            sr => \N__48239\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28647\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48757\,
            ce => \N__25153\,
            sr => \N__48241\
        );

    \current_shift_inst.un7_start_stop_0_a3_LC_4_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__48277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31028\,
            lcout => un7_start_stop_0_a3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_counter_cry_1_c_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21873\,
            in2 => \N__21556\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => un5_counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21570\,
            in2 => \_gnd_net_\,
            in3 => \N__21403\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => un5_counter_cry_1,
            carryout => un5_counter_cry_2,
            clk => \N__48867\,
            ce => 'H',
            sr => \N__48149\
        );

    \counter_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21400\,
            in2 => \_gnd_net_\,
            in3 => \N__21388\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => un5_counter_cry_2,
            carryout => un5_counter_cry_3,
            clk => \N__48867\,
            ce => 'H',
            sr => \N__48149\
        );

    \counter_4_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21385\,
            in2 => \_gnd_net_\,
            in3 => \N__21373\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => un5_counter_cry_3,
            carryout => un5_counter_cry_4,
            clk => \N__48867\,
            ce => 'H',
            sr => \N__48149\
        );

    \counter_5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21370\,
            in2 => \_gnd_net_\,
            in3 => \N__21358\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => un5_counter_cry_4,
            carryout => un5_counter_cry_5,
            clk => \N__48867\,
            ce => 'H',
            sr => \N__48149\
        );

    \counter_6_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21657\,
            in2 => \_gnd_net_\,
            in3 => \N__21643\,
            lcout => \counterZ0Z_6\,
            ltout => OPEN,
            carryin => un5_counter_cry_5,
            carryout => un5_counter_cry_6,
            clk => \N__48867\,
            ce => 'H',
            sr => \N__48149\
        );

    \counter_RNO_0_7_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21583\,
            in2 => \_gnd_net_\,
            in3 => \N__21631\,
            lcout => \counter_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => un5_counter_cry_6,
            carryout => un5_counter_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_8_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21807\,
            in2 => \_gnd_net_\,
            in3 => \N__21628\,
            lcout => \counterZ0Z_8\,
            ltout => OPEN,
            carryin => un5_counter_cry_7,
            carryout => un5_counter_cry_8,
            clk => \N__48867\,
            ce => 'H',
            sr => \N__48149\
        );

    \counter_9_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21835\,
            in2 => \_gnd_net_\,
            in3 => \N__21625\,
            lcout => \counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => un5_counter_cry_9,
            clk => \N__48861\,
            ce => 'H',
            sr => \N__48155\
        );

    \counter_RNO_0_10_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21595\,
            in2 => \_gnd_net_\,
            in3 => \N__21613\,
            lcout => \counter_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => un5_counter_cry_9,
            carryout => un5_counter_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_11_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21847\,
            in2 => \_gnd_net_\,
            in3 => \N__21610\,
            lcout => \counterZ0Z_11\,
            ltout => OPEN,
            carryin => un5_counter_cry_10,
            carryout => un5_counter_cry_11,
            clk => \N__48861\,
            ce => 'H',
            sr => \N__48155\
        );

    \counter_RNO_0_12_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21822\,
            in2 => \_gnd_net_\,
            in3 => \N__21607\,
            lcout => \counter_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI800G_7_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21594\,
            in2 => \_gnd_net_\,
            in3 => \N__21582\,
            lcout => OPEN,
            ltout => \un2_counter_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI3BSP_1_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21571\,
            in1 => \N__21548\,
            in2 => \N__21877\,
            in3 => \N__21865\,
            lcout => un2_counter_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIM6001_12_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21846\,
            in1 => \N__21834\,
            in2 => \N__21823\,
            in3 => \N__21808\,
            lcout => un2_counter_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_10khz_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__21793\,
            in1 => \N__21747\,
            in2 => \N__21691\,
            in3 => \N__21717\,
            lcout => clk_10khz_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48848\,
            ce => 'H',
            sr => \N__48178\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__35774\,
            in1 => \N__35713\,
            in2 => \N__36450\,
            in3 => \N__36655\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36658\,
            in1 => \N__36439\,
            in2 => \N__35266\,
            in3 => \N__35777\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36660\,
            in1 => \N__36441\,
            in2 => \_gnd_net_\,
            in3 => \N__36496\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36440\,
            in1 => \N__36150\,
            in2 => \_gnd_net_\,
            in3 => \N__36659\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__36656\,
            in1 => \N__35775\,
            in2 => \N__35380\,
            in3 => \N__36437\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__35773\,
            in1 => \N__35841\,
            in2 => \N__36449\,
            in3 => \N__36654\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__36657\,
            in1 => \N__35776\,
            in2 => \N__36094\,
            in3 => \N__36438\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48842\,
            ce => \N__24637\,
            sr => \N__48187\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23375\,
            in1 => \N__23498\,
            in2 => \N__23625\,
            in3 => \N__22576\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23494\,
            in1 => \N__23597\,
            in2 => \N__23392\,
            in3 => \N__22858\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23376\,
            in1 => \N__23499\,
            in2 => \N__23626\,
            in3 => \N__22822\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23495\,
            in1 => \N__23604\,
            in2 => \N__23393\,
            in3 => \N__22543\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23377\,
            in1 => \N__23500\,
            in2 => \N__23627\,
            in3 => \N__22090\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23496\,
            in1 => \N__23605\,
            in2 => \N__23394\,
            in3 => \N__22474\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23378\,
            in1 => \N__23501\,
            in2 => \N__23628\,
            in3 => \N__22441\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23497\,
            in1 => \N__23609\,
            in2 => \N__23395\,
            in3 => \N__22408\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48838\,
            ce => 'H',
            sr => \N__48195\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21886\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22000\,
            in2 => \N__22012\,
            in3 => \N__22286\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21982\,
            in2 => \N__21994\,
            in3 => \N__22554\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21964\,
            in2 => \N__21976\,
            in3 => \N__22518\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21946\,
            in2 => \N__21958\,
            in3 => \N__22485\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21925\,
            in2 => \N__21940\,
            in3 => \N__22452\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21919\,
            in2 => \N__24679\,
            in3 => \N__22419\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21913\,
            in2 => \N__24667\,
            in3 => \N__23254\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21892\,
            in2 => \N__21907\,
            in3 => \N__23230\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22069\,
            in2 => \N__22363\,
            in3 => \N__23203\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22063\,
            in2 => \N__23104\,
            in3 => \N__22764\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22737\,
            in1 => \N__22057\,
            in2 => \N__22348\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22051\,
            in2 => \N__24652\,
            in3 => \N__22710\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22045\,
            in2 => \N__23089\,
            in3 => \N__22686\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22653\,
            in1 => \N__22039\,
            in2 => \N__23119\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22623\,
            in1 => \N__23149\,
            in2 => \N__22033\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23647\,
            in1 => \N__22024\,
            in2 => \N__23071\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22018\,
            in2 => \N__22330\,
            in3 => \N__22593\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22105\,
            in2 => \N__22315\,
            in3 => \N__22875\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22839\,
            in1 => \N__22099\,
            in2 => \N__23134\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22093\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24594\,
            in1 => \N__22296\,
            in2 => \_gnd_net_\,
            in3 => \N__24541\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27967\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48803\,
            ce => \N__25134\,
            sr => \N__48219\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101010001111"
        )
    port map (
            in0 => \N__23746\,
            in1 => \N__25677\,
            in2 => \N__25558\,
            in3 => \N__25294\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48803\,
            ce => \N__25134\,
            sr => \N__48219\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__23913\,
            in1 => \_gnd_net_\,
            in2 => \N__23890\,
            in3 => \N__23937\,
            lcout => \current_shift_inst.PI_CTRL.un1_enablelt3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB4HQ_8_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24032\,
            in2 => \_gnd_net_\,
            in3 => \N__24077\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI4JA22_5_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__23690\,
            in1 => \N__23730\,
            in2 => \N__22072\,
            in3 => \N__23765\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110001"
        )
    port map (
            in0 => \N__23816\,
            in1 => \N__23844\,
            in2 => \N__22165\,
            in3 => \N__22162\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24033\,
            in1 => \N__23729\,
            in2 => \N__23694\,
            in3 => \N__23764\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23817\,
            in1 => \N__23843\,
            in2 => \N__22156\,
            in3 => \N__24078\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28450\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => \N__25135\,
            sr => \N__48226\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28012\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => \N__25135\,
            sr => \N__48226\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28147\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => \N__25135\,
            sr => \N__48226\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28801\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => \N__25135\,
            sr => \N__48226\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28060\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => \N__25135\,
            sr => \N__48226\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28369\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48785\,
            ce => \N__25135\,
            sr => \N__48226\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28723\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__25145\,
            sr => \N__48231\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24103\,
            in1 => \N__25696\,
            in2 => \N__25550\,
            in3 => \N__25336\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__25145\,
            sr => \N__48231\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28612\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__25145\,
            sr => \N__48231\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28332\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__25145\,
            sr => \N__48231\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28537\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__25145\,
            sr => \N__48231\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48776\,
            ce => \N__25145\,
            sr => \N__48231\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28293\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48767\,
            ce => \N__25178\,
            sr => \N__48234\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_5_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29032\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48758\,
            ce => \N__25194\,
            sr => \N__48237\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27343\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48751\,
            ce => \N__25179\,
            sr => \N__48240\
        );

    \pwm_generator_inst.threshold_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22384\,
            lcout => \pwm_generator_inst.thresholdZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48855\,
            ce => 'H',
            sr => \N__48139\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111110011"
        )
    port map (
            in0 => \N__29122\,
            in1 => \N__33456\,
            in2 => \N__35313\,
            in3 => \N__33633\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48849\,
            ce => 'H',
            sr => \N__48145\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24369\,
            in1 => \N__33650\,
            in2 => \_gnd_net_\,
            in3 => \N__30480\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48843\,
            ce => 'H',
            sr => \N__48150\
        );

    \pwm_generator_inst.threshold_5_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22375\,
            lcout => \pwm_generator_inst.thresholdZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48843\,
            ce => 'H',
            sr => \N__48150\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__33649\,
            in1 => \N__29209\,
            in2 => \N__35378\,
            in3 => \N__33460\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48843\,
            ce => 'H',
            sr => \N__48150\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__35986\,
            in1 => \N__35790\,
            in2 => \N__36451\,
            in3 => \N__36614\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48820\,
            ce => \N__24626\,
            sr => \N__48179\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36443\,
            in1 => \N__35889\,
            in2 => \_gnd_net_\,
            in3 => \N__36611\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48820\,
            ce => \N__24626\,
            sr => \N__48179\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__36444\,
            in1 => \N__33258\,
            in2 => \_gnd_net_\,
            in3 => \N__36612\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48820\,
            ce => \N__24626\,
            sr => \N__48179\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__36613\,
            in1 => \N__36445\,
            in2 => \_gnd_net_\,
            in3 => \N__33210\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48820\,
            ce => \N__24626\,
            sr => \N__48179\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22810\,
            in2 => \N__22300\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22561\,
            in2 => \_gnd_net_\,
            in3 => \N__22531\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23185\,
            in2 => \N__22528\,
            in3 => \N__22495\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22492\,
            in2 => \_gnd_net_\,
            in3 => \N__22462\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22459\,
            in2 => \_gnd_net_\,
            in3 => \N__22429\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22426\,
            in2 => \_gnd_net_\,
            in3 => \N__22396\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23250\,
            in2 => \_gnd_net_\,
            in3 => \N__22393\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23229\,
            in2 => \_gnd_net_\,
            in3 => \N__22390\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23199\,
            in2 => \_gnd_net_\,
            in3 => \N__22387\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22768\,
            in2 => \_gnd_net_\,
            in3 => \N__22744\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22741\,
            in2 => \_gnd_net_\,
            in3 => \N__22717\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22714\,
            in2 => \_gnd_net_\,
            in3 => \N__22690\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22687\,
            in2 => \_gnd_net_\,
            in3 => \N__22660\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22657\,
            in2 => \_gnd_net_\,
            in3 => \N__22633\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22630\,
            in2 => \_gnd_net_\,
            in3 => \N__22603\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23646\,
            in2 => \_gnd_net_\,
            in3 => \N__22600\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22597\,
            in2 => \_gnd_net_\,
            in3 => \N__22564\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22879\,
            in2 => \_gnd_net_\,
            in3 => \N__22846\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22843\,
            in2 => \_gnd_net_\,
            in3 => \N__22825\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24586\,
            in2 => \_gnd_net_\,
            in3 => \N__24542\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23438\,
            in2 => \_gnd_net_\,
            in3 => \N__23306\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24968\,
            in1 => \N__24922\,
            in2 => \N__24901\,
            in3 => \N__24821\,
            lcout => \current_shift_inst.PI_CTRL.N_47_16\,
            ltout => \current_shift_inst.PI_CTRL.N_47_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIBHHP7_18_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22912\,
            in1 => \N__22789\,
            in2 => \N__22801\,
            in3 => \N__24183\,
            lcout => \current_shift_inst.PI_CTRL.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22924\,
            in1 => \N__22774\,
            in2 => \N__26542\,
            in3 => \N__22798\,
            lcout => \current_shift_inst.PI_CTRL.N_47_21\,
            ltout => \current_shift_inst.PI_CTRL.N_47_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNITMGQ3_18_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25478\,
            in1 => \N__22783\,
            in2 => \N__22777\,
            in3 => \N__24168\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26646\,
            in1 => \N__26677\,
            in2 => \N__26613\,
            in3 => \N__26563\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26742\,
            in1 => \N__26820\,
            in2 => \N__26190\,
            in3 => \N__26783\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOU8U3_18_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24169\,
            in1 => \N__24858\,
            in2 => \N__25526\,
            in3 => \N__22890\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIE7HME_18_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__22918\,
            in1 => \N__22908\,
            in2 => \N__22894\,
            in3 => \N__26206\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1IOH6_18_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26205\,
            in1 => \N__24859\,
            in2 => \N__24179\,
            in3 => \N__22891\,
            lcout => \current_shift_inst.PI_CTRL.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24139\,
            in1 => \N__25622\,
            in2 => \N__25549\,
            in3 => \N__25293\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__25208\,
            sr => \N__48220\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__23992\,
            in1 => \N__25614\,
            in2 => \N__25547\,
            in3 => \N__25289\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__25208\,
            sr => \N__48220\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__25290\,
            in1 => \N__25509\,
            in2 => \N__25655\,
            in3 => \N__23980\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__25208\,
            sr => \N__48220\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__23947\,
            in1 => \N__25621\,
            in2 => \N__25548\,
            in3 => \N__25292\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__25208\,
            sr => \N__48220\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__25291\,
            in1 => \N__25510\,
            in2 => \N__25656\,
            in3 => \N__23971\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48768\,
            ce => \N__25208\,
            sr => \N__48220\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24115\,
            in1 => \N__25671\,
            in2 => \N__25545\,
            in3 => \N__25322\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48759\,
            ce => \N__25173\,
            sr => \N__48223\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24091\,
            in1 => \N__25672\,
            in2 => \N__25546\,
            in3 => \N__25323\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48759\,
            ce => \N__25173\,
            sr => \N__48223\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100010001"
        )
    port map (
            in0 => \N__25324\,
            in1 => \N__25499\,
            in2 => \N__25697\,
            in3 => \N__24001\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48759\,
            ce => \N__25173\,
            sr => \N__48223\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24196\,
            in1 => \N__25670\,
            in2 => \N__25544\,
            in3 => \N__25321\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48759\,
            ce => \N__25173\,
            sr => \N__48223\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28485\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48752\,
            ce => \N__25209\,
            sr => \N__48227\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28572\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48752\,
            ce => \N__25209\,
            sr => \N__48227\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28407\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48752\,
            ce => \N__25209\,
            sr => \N__48227\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24211\,
            in1 => \N__25676\,
            in2 => \N__25521\,
            in3 => \N__25325\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48752\,
            ce => \N__25209\,
            sr => \N__48227\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28996\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48752\,
            ce => \N__25209\,
            sr => \N__48227\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48746\,
            ce => \N__25195\,
            sr => \N__48232\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33781\,
            in2 => \_gnd_net_\,
            in3 => \N__29815\,
            lcout => \current_shift_inst.timer_s1.N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23038\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23029\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__30482\,
            in1 => \N__33249\,
            in2 => \N__33645\,
            in3 => \N__29671\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48850\,
            ce => 'H',
            sr => \N__48133\
        );

    \pwm_generator_inst.threshold_7_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23020\,
            lcout => \pwm_generator_inst.thresholdZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48850\,
            ce => 'H',
            sr => \N__48133\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__30483\,
            in1 => \N__35244\,
            in2 => \N__33646\,
            in3 => \N__29178\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48850\,
            ce => 'H',
            sr => \N__48133\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__29275\,
            in1 => \N__33613\,
            in2 => \N__35663\,
            in3 => \N__30481\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48850\,
            ce => 'H',
            sr => \N__48133\
        );

    \pwm_generator_inst.threshold_2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23011\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48844\,
            ce => 'H',
            sr => \N__48140\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24349\,
            in1 => \N__33651\,
            in2 => \_gnd_net_\,
            in3 => \N__30455\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48844\,
            ce => 'H',
            sr => \N__48140\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__30456\,
            in1 => \_gnd_net_\,
            in2 => \N__33655\,
            in3 => \N__24329\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48844\,
            ce => 'H',
            sr => \N__48140\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24365\,
            in1 => \N__24347\,
            in2 => \N__24331\,
            in3 => \N__26066\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.threshold_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23179\,
            lcout => \pwm_generator_inst.thresholdZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48830\,
            ce => 'H',
            sr => \N__48151\
        );

    \pwm_generator_inst.threshold_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23164\,
            lcout => \pwm_generator_inst.thresholdZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48830\,
            ce => 'H',
            sr => \N__48151\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35662\,
            in1 => \N__36398\,
            in2 => \_gnd_net_\,
            in3 => \N__36526\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48821\,
            ce => \N__24636\,
            sr => \N__48156\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__36396\,
            in1 => \N__33155\,
            in2 => \_gnd_net_\,
            in3 => \N__33130\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48821\,
            ce => \N__24636\,
            sr => \N__48156\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__33370\,
            in1 => \N__36397\,
            in2 => \_gnd_net_\,
            in3 => \N__36525\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48821\,
            ce => \N__24636\,
            sr => \N__48156\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36419\,
            in1 => \N__35931\,
            in2 => \_gnd_net_\,
            in3 => \N__36564\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48811\,
            ce => \N__24621\,
            sr => \N__48165\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36565\,
            in1 => \N__36420\,
            in2 => \_gnd_net_\,
            in3 => \N__36027\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48811\,
            ce => \N__24621\,
            sr => \N__48165\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__36566\,
            in1 => \N__36421\,
            in2 => \_gnd_net_\,
            in3 => \N__33310\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48811\,
            ce => \N__24621\,
            sr => \N__48165\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23440\,
            in1 => \N__23552\,
            in2 => \N__23344\,
            in3 => \N__23260\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48804\,
            ce => 'H',
            sr => \N__48180\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__23339\,
            in1 => \N__23442\,
            in2 => \N__23578\,
            in3 => \N__23236\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48804\,
            ce => 'H',
            sr => \N__48180\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23441\,
            in1 => \N__23556\,
            in2 => \N__23345\,
            in3 => \N__23209\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48804\,
            ce => 'H',
            sr => \N__48180\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__23551\,
            in1 => \N__23439\,
            in2 => \_gnd_net_\,
            in3 => \N__23307\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__35827\,
            in1 => \N__33634\,
            in2 => \_gnd_net_\,
            in3 => \N__30490\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48804\,
            ce => 'H',
            sr => \N__48180\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__24554\,
            in1 => \N__23340\,
            in2 => \N__23577\,
            in3 => \N__23465\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48793\,
            ce => \N__31454\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001001010"
        )
    port map (
            in0 => \N__23464\,
            in1 => \N__23550\,
            in2 => \N__23374\,
            in3 => \N__24555\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48793\,
            ce => \N__31454\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24587\,
            in2 => \_gnd_net_\,
            in3 => \N__24553\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__32896\,
            in1 => \N__32472\,
            in2 => \N__32733\,
            in3 => \N__32367\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48793\,
            ce => \N__31454\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29968\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.N_228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__23531\,
            in1 => \N__27532\,
            in2 => \N__23656\,
            in3 => \N__26110\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48786\,
            ce => 'H',
            sr => \N__48196\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__23444\,
            in1 => \N__23530\,
            in2 => \N__23346\,
            in3 => \N__23653\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48786\,
            ce => 'H',
            sr => \N__48196\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__23529\,
            in1 => \N__23443\,
            in2 => \_gnd_net_\,
            in3 => \N__23314\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101100001011"
        )
    port map (
            in0 => \N__24046\,
            in1 => \N__25252\,
            in2 => \N__25553\,
            in3 => \N__25651\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48777\,
            ce => \N__25197\,
            sr => \N__48204\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25248\,
            in1 => \N__25527\,
            in2 => \N__24130\,
            in3 => \N__25652\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48777\,
            ce => \N__25197\,
            sr => \N__48204\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101100001011"
        )
    port map (
            in0 => \N__23704\,
            in1 => \N__25250\,
            in2 => \N__25552\,
            in3 => \N__25650\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48777\,
            ce => \N__25197\,
            sr => \N__48204\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110100001101"
        )
    port map (
            in0 => \N__25251\,
            in1 => \N__23662\,
            in2 => \N__25554\,
            in3 => \N__25654\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48777\,
            ce => \N__25197\,
            sr => \N__48204\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__23959\,
            in1 => \N__25247\,
            in2 => \N__25551\,
            in3 => \N__25649\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48777\,
            ce => \N__25197\,
            sr => \N__48204\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25249\,
            in1 => \N__25528\,
            in2 => \N__23785\,
            in3 => \N__25653\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48777\,
            ce => \N__25197\,
            sr => \N__48204\
        );

    \current_shift_inst.PI_CTRL.integrator_0_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23930\,
            in2 => \N__28179\,
            in3 => \N__23862\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            clk => \N__48769\,
            ce => \N__25207\,
            sr => \N__48210\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_8_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23860\,
            in1 => \N__23912\,
            in2 => \N__28146\,
            in3 => \N__23893\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \N__48769\,
            ce => \N__25207\,
            sr => \N__48210\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23863\,
            in1 => \N__23885\,
            in2 => \N__28101\,
            in3 => \N__23866\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \N__48769\,
            ce => \N__25207\,
            sr => \N__48210\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1101011101111101"
        )
    port map (
            in0 => \N__23861\,
            in1 => \N__23842\,
            in2 => \N__28056\,
            in3 => \N__23821\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \N__48769\,
            ce => \N__25207\,
            sr => \N__48210\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23796\,
            in2 => \N__28011\,
            in3 => \N__23776\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23773\,
            in2 => \N__27963\,
            in3 => \N__23734\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23720\,
            in2 => \N__28492\,
            in3 => \N__23698\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23678\,
            in2 => \N__28449\,
            in3 => \N__24082\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24073\,
            in2 => \N__28408\,
            in3 => \N__24037\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24020\,
            in2 => \N__28368\,
            in3 => \N__23995\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26248\,
            in2 => \N__28333\,
            in3 => \N__23983\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26567\,
            in2 => \N__28294\,
            in3 => \N__23974\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26776\,
            in2 => \N__28255\,
            in3 => \N__23965\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26642\,
            in2 => \N__28219\,
            in3 => \N__23962\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26687\,
            in2 => \N__28800\,
            in3 => \N__23950\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26329\,
            in2 => \N__28761\,
            in3 => \N__23941\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26602\,
            in2 => \N__28722\,
            in3 => \N__24190\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28683\,
            in2 => \N__24825\,
            in3 => \N__24187\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24167\,
            in2 => \N__28648\,
            in3 => \N__24133\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24930\,
            in2 => \N__28611\,
            in3 => \N__24118\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24964\,
            in2 => \N__28573\,
            in3 => \N__24109\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26402\,
            in2 => \N__28536\,
            in3 => \N__24106\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24899\,
            in2 => \N__29073\,
            in3 => \N__24094\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26365\,
            in2 => \N__29031\,
            in3 => \N__24085\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26482\,
            in2 => \N__28995\,
            in3 => \N__24226\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26518\,
            in2 => \N__27344\,
            in3 => \N__24223\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27333\,
            in2 => \N__26440\,
            in3 => \N__24220\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26809\,
            in2 => \N__27345\,
            in3 => \N__24217\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27337\,
            in2 => \N__26738\,
            in3 => \N__24214\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26284\,
            in2 => \N__27346\,
            in3 => \N__24205\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27341\,
            in2 => \N__26180\,
            in3 => \N__24202\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27342\,
            in1 => \N__25401\,
            in2 => \_gnd_net_\,
            in3 => \N__24199\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.start_timer_s1_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001111110000"
        )
    port map (
            in0 => \N__24269\,
            in1 => \N__25805\,
            in2 => \N__29877\,
            in3 => \N__27928\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48740\,
            ce => \N__31432\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111001100"
        )
    port map (
            in0 => \N__27929\,
            in1 => \N__24283\,
            in2 => \N__25812\,
            in3 => \N__29822\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48740\,
            ce => \N__31432\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_RNO_0_LC_8_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24255\,
            in1 => \N__25793\,
            in2 => \N__29878\,
            in3 => \N__27927\,
            lcout => \current_shift_inst.N_199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.meas_state_0_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110101010"
        )
    port map (
            in0 => \N__27937\,
            in1 => \N__24262\,
            in2 => \N__29879\,
            in3 => \N__25794\,
            lcout => \current_shift_inst.meas_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48235\
        );

    \current_shift_inst.phase_valid_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100011111000"
        )
    port map (
            in0 => \N__25795\,
            in1 => \N__25757\,
            in2 => \N__24270\,
            in3 => \N__27936\,
            lcout => \current_shift_inst.phase_validZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48728\,
            ce => 'H',
            sr => \N__48235\
        );

    \delay_measurement_inst.hc_state_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__26006\,
            in1 => \N__25988\,
            in2 => \_gnd_net_\,
            in3 => \N__25969\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48857\,
            ce => \N__31465\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__25972\,
            in1 => \N__26008\,
            in2 => \_gnd_net_\,
            in3 => \N__25989\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48851\,
            ce => 'H',
            sr => \N__48124\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__25893\,
            in1 => \N__27273\,
            in2 => \_gnd_net_\,
            in3 => \N__30172\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_337_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30358\,
            in1 => \N__29204\,
            in2 => \N__29149\,
            in3 => \N__29226\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29528\,
            in1 => \N__29179\,
            in2 => \N__29497\,
            in3 => \N__29269\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINGQU3_9_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011101110"
        )
    port map (
            in0 => \N__29270\,
            in1 => \N__29456\,
            in2 => \N__24235\,
            in3 => \N__24232\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__24373\,
            in1 => \N__24348\,
            in2 => \N__24330\,
            in3 => \N__33115\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__33621\,
            in1 => \N__29461\,
            in2 => \N__35984\,
            in3 => \N__33445\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48831\,
            ce => 'H',
            sr => \N__48141\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110011111111"
        )
    port map (
            in0 => \N__29617\,
            in1 => \N__26068\,
            in2 => \N__33647\,
            in3 => \N__33442\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48831\,
            ce => 'H',
            sr => \N__48141\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__33411\,
            in1 => \N__33622\,
            in2 => \N__29353\,
            in3 => \N__30437\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48831\,
            ce => 'H',
            sr => \N__48141\
        );

    \pwm_generator_inst.threshold_4_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.thresholdZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48831\,
            ce => 'H',
            sr => \N__48141\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__33620\,
            in1 => \N__29496\,
            in2 => \N__36495\,
            in3 => \N__33444\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48831\,
            ce => 'H',
            sr => \N__48141\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__33443\,
            in1 => \N__29530\,
            in2 => \N__35423\,
            in3 => \N__33626\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48831\,
            ce => 'H',
            sr => \N__48141\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001001100"
        )
    port map (
            in0 => \N__35658\,
            in1 => \N__24295\,
            in2 => \N__26050\,
            in3 => \N__24517\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto5_3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35370\,
            in1 => \N__35691\,
            in2 => \N__36086\,
            in3 => \N__35837\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto5Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto6_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__36129\,
            in1 => \N__35315\,
            in2 => \N__24286\,
            in3 => \N__35254\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlt8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto9_0_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__33365\,
            in1 => \N__35967\,
            in2 => \N__24520\,
            in3 => \N__26074\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlt15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24493\,
            in2 => \N__24511\,
            in3 => \N__27660\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27605\,
            in1 => \N__24478\,
            in2 => \N__24487\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24457\,
            in2 => \N__24472\,
            in3 => \N__27642\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24442\,
            in2 => \N__24451\,
            in3 => \N__27584\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24424\,
            in2 => \N__24436\,
            in3 => \N__27623\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24403\,
            in2 => \N__24418\,
            in3 => \N__27719\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24379\,
            in2 => \N__24397\,
            in3 => \N__27737\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24754\,
            in2 => \N__24772\,
            in3 => \N__27755\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24730\,
            in2 => \N__24748\,
            in3 => \N__27774\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24706\,
            in2 => \N__24724\,
            in3 => \N__27792\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24700\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48805\,
            ce => 'H',
            sr => \N__48157\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__35323\,
            in1 => \N__35769\,
            in2 => \N__36442\,
            in3 => \N__36561\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48794\,
            ce => \N__24622\,
            sr => \N__48166\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36563\,
            in1 => \N__36418\,
            in2 => \_gnd_net_\,
            in3 => \N__35424\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48794\,
            ce => \N__24622\,
            sr => \N__48166\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36562\,
            in1 => \N__36417\,
            in2 => \_gnd_net_\,
            in3 => \N__33407\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48794\,
            ce => \N__24622\,
            sr => \N__48166\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__29970\,
            in1 => \N__24595\,
            in2 => \N__24565\,
            in3 => \N__24556\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48778\,
            ce => 'H',
            sr => \N__48188\
        );

    \phase_controller_inst1.state_2_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__29969\,
            in1 => \N__39583\,
            in2 => \N__29936\,
            in3 => \N__26139\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48778\,
            ce => 'H',
            sr => \N__48188\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24973\,
            in1 => \N__24923\,
            in2 => \N__24900\,
            in3 => \N__24811\,
            lcout => \current_shift_inst.PI_CTRL.N_46_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39643\,
            in2 => \_gnd_net_\,
            in3 => \N__39549\,
            lcout => \phase_controller_inst1.N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__25657\,
            in1 => \N__24844\,
            in2 => \N__25522\,
            in3 => \N__25326\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48760\,
            ce => \N__25210\,
            sr => \N__48205\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25327\,
            in1 => \N__25466\,
            in2 => \N__24838\,
            in3 => \N__25658\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48760\,
            ce => \N__25210\,
            sr => \N__48205\
        );

    \current_shift_inst.start_timer_phase_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100101010"
        )
    port map (
            in0 => \N__31784\,
            in1 => \N__25813\,
            in2 => \N__25765\,
            in3 => \N__27915\,
            lcout => \current_shift_inst.start_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48753\,
            ce => \N__31444\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24790\,
            in1 => \N__25698\,
            in2 => \N__25476\,
            in3 => \N__25328\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48747\,
            ce => \N__25174\,
            sr => \N__48215\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000001100"
        )
    port map (
            in0 => \N__25330\,
            in1 => \N__25421\,
            in2 => \N__25708\,
            in3 => \N__24784\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48747\,
            ce => \N__25174\,
            sr => \N__48215\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__24778\,
            in1 => \N__25699\,
            in2 => \N__25477\,
            in3 => \N__25329\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48747\,
            ce => \N__25174\,
            sr => \N__48215\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__25706\,
            in1 => \N__25738\,
            in2 => \N__25474\,
            in3 => \N__25334\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48741\,
            ce => \N__25196\,
            sr => \N__48221\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011101100"
        )
    port map (
            in0 => \N__25332\,
            in1 => \N__25410\,
            in2 => \N__25732\,
            in3 => \N__25704\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48741\,
            ce => \N__25196\,
            sr => \N__48221\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100100011111000"
        )
    port map (
            in0 => \N__25335\,
            in1 => \N__25723\,
            in2 => \N__25475\,
            in3 => \N__25707\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48741\,
            ce => \N__25196\,
            sr => \N__48221\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011000100"
        )
    port map (
            in0 => \N__25705\,
            in1 => \N__25417\,
            in2 => \N__25717\,
            in3 => \N__25333\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48741\,
            ce => \N__25196\,
            sr => \N__48221\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110011010000"
        )
    port map (
            in0 => \N__25703\,
            in1 => \N__25564\,
            in2 => \N__25473\,
            in3 => \N__25331\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48741\,
            ce => \N__25196\,
            sr => \N__48221\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILORI_11_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40419\,
            in2 => \_gnd_net_\,
            in3 => \N__34357\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILORI_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJDBL1_10_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40564\,
            in1 => \N__40503\,
            in2 => \N__34444\,
            in3 => \N__34401\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJDBL1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1PG21_9_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40563\,
            in2 => \_gnd_net_\,
            in3 => \N__34440\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1PG21_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR0UI_13_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40265\,
            in2 => \_gnd_net_\,
            in3 => \N__34275\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR0UI_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI53NU1_6_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \N__33916\,
            in1 => \N__39930\,
            in2 => \N__40701\,
            in3 => \N__34522\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI53NU1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHVAV_6_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__39929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33915\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHVAV_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIK3CV_7_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__40697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34521\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIK3CV_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIER9V_5_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39990\,
            in2 => \_gnd_net_\,
            in3 => \N__33960\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIER9V_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJ3381_21_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__34600\,
            in1 => \N__40764\,
            in2 => \N__34642\,
            in3 => \N__41721\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJ3381_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync0_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45684\,
            lcout => \current_shift_inst.S3_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32509\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_phase_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111000000"
        )
    port map (
            in0 => \N__27930\,
            in1 => \N__25801\,
            in2 => \N__25761\,
            in3 => \N__31750\,
            lcout => \current_shift_inst.stop_timer_phaseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48721\,
            ce => \N__31412\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100001011000"
        )
    port map (
            in0 => \N__32851\,
            in1 => \N__32731\,
            in2 => \N__32596\,
            in3 => \N__32360\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48721\,
            ce => \N__31412\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_rise_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25840\,
            in2 => \_gnd_net_\,
            in3 => \N__25848\,
            lcout => \current_shift_inst.S3_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync1_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25858\,
            lcout => \current_shift_inst.S3_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S3_sync_prev_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25849\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S3_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48276\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_10_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37966\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_hc_sig_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25970\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48845\,
            ce => 'H',
            sr => \N__48101\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_3_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25944\,
            in2 => \_gnd_net_\,
            in3 => \N__25917\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25881\,
            in1 => \N__25905\,
            in2 => \N__25822\,
            in3 => \N__25819\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_26_2_4_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25869\,
            in1 => \N__27231\,
            in2 => \N__25933\,
            in3 => \N__27243\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_26_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__26007\,
            in1 => \N__25990\,
            in2 => \N__48280\,
            in3 => \N__25971\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__25945\,
            in1 => \N__33558\,
            in2 => \_gnd_net_\,
            in3 => \N__30425\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30427\,
            in1 => \N__25932\,
            in2 => \_gnd_net_\,
            in3 => \N__33561\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__25918\,
            in1 => \N__33557\,
            in2 => \_gnd_net_\,
            in3 => \N__30424\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__30428\,
            in1 => \N__33559\,
            in2 => \N__36139\,
            in3 => \N__29148\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__25906\,
            in1 => \N__33555\,
            in2 => \_gnd_net_\,
            in3 => \N__30422\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__27274\,
            in1 => \N__25894\,
            in2 => \_gnd_net_\,
            in3 => \N__30173\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__25882\,
            in1 => \N__33556\,
            in2 => \_gnd_net_\,
            in3 => \N__30423\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30426\,
            in1 => \N__25870\,
            in2 => \_gnd_net_\,
            in3 => \N__33560\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48832\,
            ce => 'H',
            sr => \N__48117\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ0JH1_6_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29495\,
            in1 => \N__29529\,
            in2 => \N__29121\,
            in3 => \N__29271\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52G18_14_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000100"
        )
    port map (
            in0 => \N__26017\,
            in1 => \N__27481\,
            in2 => \N__26035\,
            in3 => \N__26032\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_0_31_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__27378\,
            in1 => \N__27452\,
            in2 => \N__26026\,
            in3 => \N__29721\,
            lcout => \delay_measurement_inst.delay_hc_reg3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5483B_31_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__27453\,
            in1 => \N__27379\,
            in2 => \N__29725\,
            in3 => \N__26023\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto31_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29379\,
            in1 => \N__29415\,
            in2 => \N__29352\,
            in3 => \N__29307\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOHNN2_6_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__27409\,
            in1 => \N__29457\,
            in2 => \N__26011\,
            in3 => \N__29117\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__33544\,
            in1 => \N__29227\,
            in2 => \N__35709\,
            in3 => \N__33441\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48813\,
            ce => 'H',
            sr => \N__48128\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__30419\,
            in1 => \N__29383\,
            in2 => \N__33602\,
            in3 => \N__35888\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48813\,
            ce => 'H',
            sr => \N__48128\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__30421\,
            in1 => \N__33208\,
            in2 => \N__33604\,
            in3 => \N__29644\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48813\,
            ce => 'H',
            sr => \N__48128\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__35930\,
            in1 => \N__33545\,
            in2 => \N__29419\,
            in3 => \N__30418\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48813\,
            ce => 'H',
            sr => \N__48128\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__30420\,
            in1 => \N__36018\,
            in2 => \N__33603\,
            in3 => \N__29311\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48813\,
            ce => 'H',
            sr => \N__48128\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_3_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33393\,
            in1 => \N__35868\,
            in2 => \N__36019\,
            in3 => \N__35910\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto13_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto13_3_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__36477\,
            in1 => \N__35403\,
            in2 => \N__26077\,
            in3 => \N__35966\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__33254\,
            in1 => \N__26067\,
            in2 => \N__33204\,
            in3 => \N__33307\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto19Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36020\,
            in1 => \N__35664\,
            in2 => \N__33308\,
            in3 => \N__33369\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36490\,
            in1 => \N__35416\,
            in2 => \N__36149\,
            in3 => \N__35923\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33253\,
            in1 => \N__33406\,
            in2 => \N__33209\,
            in3 => \N__35881\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27697\,
            in1 => \N__27661\,
            in2 => \_gnd_net_\,
            in3 => \N__26041\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_12_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27691\,
            in1 => \N__27607\,
            in2 => \_gnd_net_\,
            in3 => \N__26038\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27698\,
            in1 => \N__27643\,
            in2 => \_gnd_net_\,
            in3 => \N__26101\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_3_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27692\,
            in1 => \N__27586\,
            in2 => \_gnd_net_\,
            in3 => \N__26098\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_4_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27699\,
            in1 => \N__27625\,
            in2 => \_gnd_net_\,
            in3 => \N__26095\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_5_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27693\,
            in1 => \N__27720\,
            in2 => \_gnd_net_\,
            in3 => \N__26092\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_6_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27700\,
            in1 => \N__27738\,
            in2 => \_gnd_net_\,
            in3 => \N__26089\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_7_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27694\,
            in1 => \N__27757\,
            in2 => \_gnd_net_\,
            in3 => \N__26086\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__48788\,
            ce => 'H',
            sr => \N__48146\
        );

    \pwm_generator_inst.counter_8_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27696\,
            in1 => \N__27775\,
            in2 => \_gnd_net_\,
            in3 => \N__26083\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_10_13_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__48780\,
            ce => 'H',
            sr => \N__48152\
        );

    \pwm_generator_inst.counter_9_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__27793\,
            in1 => \N__27695\,
            in2 => \_gnd_net_\,
            in3 => \N__26080\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48780\,
            ce => 'H',
            sr => \N__48152\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31021\,
            in2 => \_gnd_net_\,
            in3 => \N__27526\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.N_232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__39584\,
            in1 => \N__26143\,
            in2 => \N__26146\,
            in3 => \N__27552\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48771\,
            ce => 'H',
            sr => \N__48158\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI190J_15_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__41190\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34866\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI190J_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39579\,
            in2 => \_gnd_net_\,
            in3 => \N__26138\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIIKQI_10_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40504\,
            in2 => \_gnd_net_\,
            in3 => \N__34400\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIIKQI_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPB581_22_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__34554\,
            in1 => \N__41728\,
            in2 => \N__41661\,
            in3 => \N__34596\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPB581_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDR081_20_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40843\,
            in1 => \N__40770\,
            in2 => \N__34686\,
            in3 => \N__34628\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDR081_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIH6661_17_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__41047\,
            in1 => \N__34749\,
            in2 => \N__34801\,
            in3 => \N__40984\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIH6661_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOV0K_21_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40771\,
            in2 => \_gnd_net_\,
            in3 => \N__34627\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOV0K_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5M161_15_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__41191\,
            in1 => \N__34834\,
            in2 => \N__34873\,
            in3 => \N__41111\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5M161_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__32626\,
            in1 => \N__32852\,
            in2 => \_gnd_net_\,
            in3 => \N__32499\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIR32K_22_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41727\,
            in2 => \_gnd_net_\,
            in3 => \N__34595\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIR32K_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26691\,
            in1 => \N__26641\,
            in2 => \N__26617\,
            in3 => \N__26575\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIP5T51_13_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__34276\,
            in1 => \N__40194\,
            in2 => \N__40276\,
            in3 => \N__34232\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP5T51_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26526\,
            in1 => \N__26491\,
            in2 => \N__26454\,
            in3 => \N__26406\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_1_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7OAK_29_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41247\,
            in2 => \_gnd_net_\,
            in3 => \N__34959\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7OAK_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26525\,
            in1 => \N__26489\,
            in2 => \N__26453\,
            in3 => \N__26401\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26377\,
            in1 => \N__26336\,
            in2 => \N__26302\,
            in3 => \N__26255\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA53P2_0_10_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26221\,
            in1 => \N__26215\,
            in2 => \N__26209\,
            in3 => \N__26704\,
            lcout => \current_shift_inst.PI_CTRL.N_46_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26176\,
            in1 => \N__26821\,
            in2 => \N__26785\,
            in3 => \N__26728\,
            lcout => \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNILRVJ_20_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40842\,
            in2 => \_gnd_net_\,
            in3 => \N__34685\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNILRVJ_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__37362\,
            in1 => \N__40058\,
            in2 => \_gnd_net_\,
            in3 => \N__34001\,
            lcout => \current_shift_inst.un38_control_input_0_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIOSSI_12_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40342\,
            in2 => \_gnd_net_\,
            in3 => \N__34312\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIOSSI_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_0_13_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38884\,
            in2 => \_gnd_net_\,
            in3 => \N__36822\,
            lcout => \phase_controller_inst1.stoper_tr.N_21\,
            ltout => \phase_controller_inst1.stoper_tr.N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26698\,
            in3 => \N__45154\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU4VI_14_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40195\,
            in2 => \_gnd_net_\,
            in3 => \N__34234\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU4VI_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIE6961_18_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40983\,
            in1 => \N__40905\,
            in2 => \N__34759\,
            in3 => \N__34723\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIE6961_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAL3J_18_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40982\,
            in2 => \_gnd_net_\,
            in3 => \N__34755\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAL3J_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIO0U12_8_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__34486\,
            in1 => \N__40562\,
            in2 => \N__40636\,
            in3 => \N__34439\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIO0U12_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_RNO_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__34108\,
            in1 => \N__37444\,
            in2 => \_gnd_net_\,
            in3 => \N__37329\,
            lcout => \current_shift_inst.un38_control_input_0_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_0_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40059\,
            in2 => \_gnd_net_\,
            in3 => \N__34002\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNO_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40060\,
            in1 => \N__39989\,
            in2 => \N__34006\,
            in3 => \N__33953\,
            lcout => \current_shift_inst.un38_control_input_0_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_RNO_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110010011100"
        )
    port map (
            in0 => \N__37330\,
            in1 => \N__37294\,
            in2 => \N__37450\,
            in3 => \N__34069\,
            lcout => \current_shift_inst.un38_control_input_0_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CRY_0_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37448\,
            in2 => \N__37449\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_0_c_inv_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26857\,
            in2 => \N__34171\,
            in3 => \N__34893\,
            lcout => \current_shift_inst.z_i_0_31\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0_c_THRU_CO\,
            carryout => \current_shift_inst.un38_control_input_0_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_1_c_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34107\,
            in2 => \N__26851\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_0\,
            carryout => \current_shift_inst.un38_control_input_0_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_2_c_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34065\,
            in2 => \N__26839\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_1\,
            carryout => \current_shift_inst.un38_control_input_0_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34033\,
            in2 => \N__26830\,
            in3 => \N__37465\,
            lcout => \current_shift_inst.un38_control_input_0_cry_3_c_invZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_2\,
            carryout => \current_shift_inst.un38_control_input_0_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_4_c_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26977\,
            in2 => \N__37363\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_3\,
            carryout => \current_shift_inst.un38_control_input_0_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26968\,
            in2 => \N__26959\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_4\,
            carryout => \current_shift_inst.un38_control_input_0_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_5_c_RNI7HN13_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30079\,
            in2 => \N__26947\,
            in3 => \N__26938\,
            lcout => \current_shift_inst.control_input_1_axb_0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_5\,
            carryout => \current_shift_inst.un38_control_input_0_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_6_c_RNIHVR13_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26935\,
            in2 => \N__26929\,
            in3 => \N__26917\,
            lcout => \current_shift_inst.control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_7_c_RNIRD023_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31621\,
            in2 => \N__26914\,
            in3 => \N__26905\,
            lcout => \current_shift_inst.control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_7\,
            carryout => \current_shift_inst.un38_control_input_0_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_8_c_RNIC9753_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26902\,
            in2 => \N__31375\,
            in3 => \N__26893\,
            lcout => \current_shift_inst.control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_8\,
            carryout => \current_shift_inst.un38_control_input_0_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_9_c_RNII9PR2_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26890\,
            in2 => \N__26884\,
            in3 => \N__26875\,
            lcout => \current_shift_inst.control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_9\,
            carryout => \current_shift_inst.un38_control_input_0_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_10_c_RNIV96V1_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27817\,
            in2 => \N__26872\,
            in3 => \N__26860\,
            lcout => \current_shift_inst.control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_10\,
            carryout => \current_shift_inst.un38_control_input_0_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_11_c_RNI9OAV1_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31588\,
            in2 => \N__27112\,
            in3 => \N__27103\,
            lcout => \current_shift_inst.control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_11\,
            carryout => \current_shift_inst.un38_control_input_0_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_12_c_RNIJ6FV1_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31555\,
            in2 => \N__27100\,
            in3 => \N__27088\,
            lcout => \current_shift_inst.control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_12\,
            carryout => \current_shift_inst.un38_control_input_0_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_13_c_RNITKJV1_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27085\,
            in2 => \N__27079\,
            in3 => \N__27067\,
            lcout => \current_shift_inst.control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_13\,
            carryout => \current_shift_inst.un38_control_input_0_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_14_c_RNI73OV1_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31540\,
            in2 => \N__27064\,
            in3 => \N__27052\,
            lcout => \current_shift_inst.control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_15_c_RNIHHSV1_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27049\,
            in2 => \N__27037\,
            in3 => \N__27025\,
            lcout => \current_shift_inst.control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_15\,
            carryout => \current_shift_inst.un38_control_input_0_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_16_c_RNIRV002_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31510\,
            in2 => \N__31483\,
            in3 => \N__27022\,
            lcout => \current_shift_inst.control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_16\,
            carryout => \current_shift_inst.un38_control_input_0_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_17_c_RNI5E502_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27019\,
            in2 => \N__34189\,
            in3 => \N__27010\,
            lcout => \current_shift_inst.control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_17\,
            carryout => \current_shift_inst.un38_control_input_0_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_18_c_RNI6KA02_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27007\,
            in2 => \N__26998\,
            in3 => \N__26983\,
            lcout => \current_shift_inst.control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_18\,
            carryout => \current_shift_inst.un38_control_input_0_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_19_c_RNICO912_LC_10_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31525\,
            in2 => \N__31609\,
            in3 => \N__26980\,
            lcout => \current_shift_inst.control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_19\,
            carryout => \current_shift_inst.un38_control_input_0_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_20_c_RNI92P32_LC_10_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27208\,
            in2 => \N__27199\,
            in3 => \N__27187\,
            lcout => \current_shift_inst.control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_20\,
            carryout => \current_shift_inst.un38_control_input_0_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_21_c_RNIJGT32_LC_10_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27184\,
            in2 => \N__27178\,
            in3 => \N__27166\,
            lcout => \current_shift_inst.control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_21\,
            carryout => \current_shift_inst.un38_control_input_0_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_22_c_RNITU142_LC_10_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27163\,
            in2 => \N__27148\,
            in3 => \N__27130\,
            lcout => \current_shift_inst.control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \bfn_10_24_0_\,
            carryout => \current_shift_inst.un38_control_input_0_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_23_c_RNI7D642_LC_10_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28837\,
            in2 => \N__31573\,
            in3 => \N__27127\,
            lcout => \current_shift_inst.control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_23\,
            carryout => \current_shift_inst.un38_control_input_0_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_24_c_RNIHRA42_LC_10_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31666\,
            in2 => \N__28831\,
            in3 => \N__27124\,
            lcout => \current_shift_inst.control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_24\,
            carryout => \current_shift_inst.un38_control_input_0_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_25_c_RNIR9F42_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31651\,
            in2 => \N__28822\,
            in3 => \N__27121\,
            lcout => \current_shift_inst.control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_25\,
            carryout => \current_shift_inst.un38_control_input_0_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_26_c_RNI5OJ42_LC_10_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31807\,
            in2 => \N__31720\,
            in3 => \N__27118\,
            lcout => \current_shift_inst.control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_26\,
            carryout => \current_shift_inst.un38_control_input_0_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_27_c_RNIF6O42_LC_10_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31636\,
            in2 => \N__31699\,
            in3 => \N__27115\,
            lcout => \current_shift_inst.control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_27\,
            carryout => \current_shift_inst.un38_control_input_0_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_28_c_RNIGCT42_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31681\,
            in2 => \N__27832\,
            in3 => \N__27355\,
            lcout => \current_shift_inst.control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_28\,
            carryout => \current_shift_inst.un38_control_input_0_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_0_cry_29_c_RNIMGS52_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28843\,
            in2 => \N__28866\,
            in3 => \N__27352\,
            lcout => \current_shift_inst.control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_0_cry_29\,
            carryout => \current_shift_inst.un38_control_input_0_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_25_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31495\,
            in2 => \N__28879\,
            in3 => \N__27349\,
            lcout => \current_shift_inst.control_inputZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48704\,
            ce => \N__28963\,
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27272\,
            in2 => \_gnd_net_\,
            in3 => \N__30174\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_336_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__27244\,
            in1 => \N__33586\,
            in2 => \_gnd_net_\,
            in3 => \N__30467\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48833\,
            ce => 'H',
            sr => \N__48102\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__30468\,
            in1 => \_gnd_net_\,
            in2 => \N__33627\,
            in3 => \N__27232\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48833\,
            ce => 'H',
            sr => \N__48102\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27220\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJD01_11_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29348\,
            in1 => \N__29372\,
            in2 => \N__30519\,
            in3 => \N__29268\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29475\,
            in2 => \_gnd_net_\,
            in3 => \N__29511\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_10_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27403\,
            in1 => \N__27394\,
            in2 => \N__27397\,
            in3 => \N__27385\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOKRB1_10_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__29616\,
            in1 => \N__30356\,
            in2 => \N__29208\,
            in3 => \N__29405\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29637\,
            in2 => \_gnd_net_\,
            in3 => \N__29664\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4UNN2_4_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__27475\,
            in1 => \N__29171\,
            in2 => \N__27388\,
            in3 => \N__29144\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP8VO1_20_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__29569\,
            in1 => \N__27468\,
            in2 => \N__29557\,
            in3 => \N__29587\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29553\,
            in2 => \_gnd_net_\,
            in3 => \N__29568\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1LC84_14_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__30515\,
            in1 => \N__27370\,
            in2 => \N__27493\,
            in3 => \N__29267\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1lt30_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOVQ9D_14_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27364\,
            in1 => \N__27457\,
            in2 => \N__27358\,
            in3 => \N__27499\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINN412_20_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__29586\,
            in1 => \N__27469\,
            in2 => \N__29720\,
            in3 => \N__27505\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29636\,
            in1 => \N__29663\,
            in2 => \N__29615\,
            in3 => \N__29990\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30511\,
            in2 => \N__27484\,
            in3 => \N__29266\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2VRB1_13_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29438\,
            in1 => \N__29100\,
            in2 => \N__29306\,
            in3 => \N__29991\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29788\,
            in1 => \N__29797\,
            in2 => \N__29779\,
            in3 => \N__29539\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29749\,
            in1 => \N__29758\,
            in2 => \N__29740\,
            in3 => \N__29767\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_13_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27433\,
            in1 => \N__27427\,
            in2 => \N__27421\,
            in3 => \N__27799\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33159\,
            in2 => \N__27412\,
            in3 => \N__33125\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlt31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35314\,
            in1 => \N__35985\,
            in2 => \_gnd_net_\,
            in3 => \N__35255\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__36087\,
            in1 => \N__35379\,
            in2 => \N__27802\,
            in3 => \N__35704\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27791\,
            in1 => \N__27773\,
            in2 => \_gnd_net_\,
            in3 => \N__27756\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27739\,
            in1 => \N__27721\,
            in2 => \N__27703\,
            in3 => \N__27568\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27659\,
            in2 => \_gnd_net_\,
            in3 => \N__27641\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__27624\,
            in1 => \N__27606\,
            in2 => \N__27589\,
            in3 => \N__27585\,
            lcout => \pwm_generator_inst.un1_counterlt9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27562\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48761\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__31792\,
            in1 => \N__31831\,
            in2 => \_gnd_net_\,
            in3 => \N__31762\,
            lcout => \current_shift_inst.timer_phase.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48755\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.start_timer_tr_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__27528\,
            in1 => \N__27853\,
            in2 => \N__32684\,
            in3 => \N__27553\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48755\,
            ce => 'H',
            sr => \N__48159\
        );

    \phase_controller_inst1.state_4_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30984\,
            in2 => \_gnd_net_\,
            in3 => \N__27527\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48755\,
            ce => 'H',
            sr => \N__48159\
        );

    \current_shift_inst.S1_rise_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27838\,
            in2 => \_gnd_net_\,
            in3 => \N__27846\,
            lcout => \current_shift_inst.S1_riseZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync0_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30030\,
            lcout => \current_shift_inst.S1_syncZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync1_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27859\,
            lcout => \current_shift_inst.S1_syncZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39666\,
            in2 => \_gnd_net_\,
            in3 => \N__29903\,
            lcout => \phase_controller_inst1.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.S1_sync_prev_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.S1_sync_prevZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48749\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__29904\,
            in1 => \N__39635\,
            in2 => \N__39683\,
            in3 => \N__39545\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48743\,
            ce => 'H',
            sr => \N__48181\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__49126\,
            in1 => \N__47179\,
            in2 => \_gnd_net_\,
            in3 => \N__46240\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48736\,
            ce => \N__46354\,
            sr => \N__48189\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIKKJ81_29_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__41336\,
            in1 => \N__34960\,
            in2 => \N__35002\,
            in3 => \N__41248\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIKKJ81_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7DM51_10_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40502\,
            in1 => \N__34355\,
            in2 => \N__34402\,
            in3 => \N__40412\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7DM51_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39814\,
            in1 => \N__39763\,
            in2 => \N__39736\,
            in3 => \N__45253\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__45153\,
            in1 => \N__45057\,
            in2 => \_gnd_net_\,
            in3 => \N__44994\,
            lcout => \phase_controller_inst1.stoper_tr.N_20_li\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_0_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28189\,
            in2 => \N__30094\,
            in3 => \N__30093\,
            lcout => \current_shift_inst.control_inputZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \current_shift_inst.control_input_1_cry_0\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28156\,
            in2 => \_gnd_net_\,
            in3 => \N__28117\,
            lcout => \current_shift_inst.control_inputZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_0\,
            carryout => \current_shift_inst.control_input_1_cry_1\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_2_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28114\,
            in2 => \_gnd_net_\,
            in3 => \N__28072\,
            lcout => \current_shift_inst.control_inputZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_1\,
            carryout => \current_shift_inst.control_input_1_cry_2\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_3_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28069\,
            in2 => \_gnd_net_\,
            in3 => \N__28027\,
            lcout => \current_shift_inst.control_inputZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_2\,
            carryout => \current_shift_inst.control_input_1_cry_3\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_4_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28024\,
            in3 => \N__27982\,
            lcout => \current_shift_inst.control_inputZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_3\,
            carryout => \current_shift_inst.control_input_1_cry_4\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_5_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27979\,
            in3 => \N__27940\,
            lcout => \current_shift_inst.control_inputZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_4\,
            carryout => \current_shift_inst.control_input_1_cry_5\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_6_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28504\,
            in3 => \N__28465\,
            lcout => \current_shift_inst.control_inputZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_5\,
            carryout => \current_shift_inst.control_input_1_cry_6\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_7_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28462\,
            in3 => \N__28420\,
            lcout => \current_shift_inst.control_inputZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_6\,
            carryout => \current_shift_inst.control_input_1_cry_7\,
            clk => \N__48723\,
            ce => \N__28950\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_8_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28417\,
            in3 => \N__28381\,
            lcout => \current_shift_inst.control_inputZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_21_0_\,
            carryout => \current_shift_inst.control_input_1_cry_8\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_9_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28378\,
            in2 => \_gnd_net_\,
            in3 => \N__28345\,
            lcout => \current_shift_inst.control_inputZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_8\,
            carryout => \current_shift_inst.control_input_1_cry_9\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_10_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28342\,
            in2 => \_gnd_net_\,
            in3 => \N__28306\,
            lcout => \current_shift_inst.control_inputZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_9\,
            carryout => \current_shift_inst.control_input_1_cry_10\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_11_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28303\,
            in2 => \_gnd_net_\,
            in3 => \N__28267\,
            lcout => \current_shift_inst.control_inputZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_10\,
            carryout => \current_shift_inst.control_input_1_cry_11\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_12_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28264\,
            in2 => \_gnd_net_\,
            in3 => \N__28234\,
            lcout => \current_shift_inst.control_inputZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_11\,
            carryout => \current_shift_inst.control_input_1_cry_12\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_13_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28231\,
            in3 => \N__28192\,
            lcout => \current_shift_inst.control_inputZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_12\,
            carryout => \current_shift_inst.control_input_1_cry_13\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_14_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28813\,
            in3 => \N__28777\,
            lcout => \current_shift_inst.control_inputZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_13\,
            carryout => \current_shift_inst.control_input_1_cry_14\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_15_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28774\,
            in3 => \N__28732\,
            lcout => \current_shift_inst.control_inputZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_14\,
            carryout => \current_shift_inst.control_input_1_cry_15\,
            clk => \N__48716\,
            ce => \N__28964\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_16_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28729\,
            in2 => \_gnd_net_\,
            in3 => \N__28696\,
            lcout => \current_shift_inst.control_inputZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \current_shift_inst.control_input_1_cry_16\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_17_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28693\,
            in2 => \_gnd_net_\,
            in3 => \N__28660\,
            lcout => \current_shift_inst.control_inputZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_16\,
            carryout => \current_shift_inst.control_input_1_cry_17\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_18_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28657\,
            in2 => \_gnd_net_\,
            in3 => \N__28624\,
            lcout => \current_shift_inst.control_inputZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_17\,
            carryout => \current_shift_inst.control_input_1_cry_18\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_19_LC_11_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28621\,
            in2 => \_gnd_net_\,
            in3 => \N__28588\,
            lcout => \current_shift_inst.control_inputZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_18\,
            carryout => \current_shift_inst.control_input_1_cry_19\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_20_LC_11_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28585\,
            in3 => \N__28552\,
            lcout => \current_shift_inst.control_inputZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_19\,
            carryout => \current_shift_inst.control_input_1_cry_20\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_21_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28549\,
            in3 => \N__28507\,
            lcout => \current_shift_inst.control_inputZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_20\,
            carryout => \current_shift_inst.control_input_1_cry_21\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_22_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29086\,
            in3 => \N__29047\,
            lcout => \current_shift_inst.control_inputZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_21\,
            carryout => \current_shift_inst.control_input_1_cry_22\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_23_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29044\,
            in3 => \N__29005\,
            lcout => \current_shift_inst.control_inputZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_1_cry_22\,
            carryout => \current_shift_inst.control_input_1_cry_23\,
            clk => \N__48710\,
            ce => \N__28965\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_24_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29002\,
            in2 => \_gnd_net_\,
            in3 => \N__28972\,
            lcout => \current_shift_inst.control_inputZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \current_shift_inst.control_input_1_cry_24\,
            clk => \N__48707\,
            ce => \N__28969\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_1_cry_24_THRU_LUT4_0_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28882\,
            lcout => \current_shift_inst.control_input_1_cry_24_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQF91_30_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__28867\,
            in1 => \N__41886\,
            in2 => \_gnd_net_\,
            in3 => \N__34927\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQF91_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVJ781_23_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111000011"
        )
    port map (
            in0 => \N__34558\,
            in1 => \N__41579\,
            in2 => \N__35131\,
            in3 => \N__41654\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVJ781_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI1C4K_24_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__41580\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35130\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI1C4K_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4G5K_25_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41520\,
            in2 => \_gnd_net_\,
            in3 => \N__35095\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4G5K_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__32686\,
            in1 => \N__32895\,
            in2 => \N__30199\,
            in3 => \N__32569\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48702\,
            ce => 'H',
            sr => \N__48228\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_11_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__32685\,
            in1 => \N__32894\,
            in2 => \_gnd_net_\,
            in3 => \N__32568\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_11_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__39631\,
            in1 => \N__32406\,
            in2 => \N__29230\,
            in3 => \N__32368\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48702\,
            ce => 'H',
            sr => \N__48228\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30337\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48822\,
            ce => \N__29691\,
            sr => \N__48095\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30316\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48822\,
            ce => \N__29691\,
            sr => \N__48095\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30336\,
            in2 => \N__30294\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30315\,
            in2 => \N__30270\,
            in3 => \N__29152\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30245\,
            in2 => \N__30295\,
            in3 => \N__29125\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30227\,
            in2 => \N__30271\,
            in3 => \N__29089\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30246\,
            in2 => \N__30726\,
            in3 => \N__29500\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30228\,
            in2 => \N__30702\,
            in3 => \N__29464\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30679\,
            in2 => \N__30727\,
            in3 => \N__29422\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30655\,
            in2 => \N__30703\,
            in3 => \N__29386\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__48812\,
            ce => \N__29692\,
            sr => \N__48103\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30678\,
            in2 => \N__30630\,
            in3 => \N__29356\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30654\,
            in2 => \N__30606\,
            in3 => \N__29314\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30581\,
            in2 => \N__30631\,
            in3 => \N__29281\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30563\,
            in2 => \N__30607\,
            in3 => \N__29278\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30582\,
            in2 => \N__30546\,
            in3 => \N__29233\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30564\,
            in2 => \N__30906\,
            in3 => \N__29674\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30883\,
            in2 => \N__30547\,
            in3 => \N__29647\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30859\,
            in2 => \N__30907\,
            in3 => \N__29620\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__48806\,
            ce => \N__29693\,
            sr => \N__48109\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30882\,
            in2 => \N__30834\,
            in3 => \N__29590\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30858\,
            in2 => \N__30810\,
            in3 => \N__29572\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30785\,
            in2 => \N__30835\,
            in3 => \N__29560\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30767\,
            in2 => \N__30811\,
            in3 => \N__29542\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30786\,
            in2 => \N__30750\,
            in3 => \N__29533\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30768\,
            in2 => \N__31356\,
            in3 => \N__29791\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31333\,
            in2 => \N__30751\,
            in3 => \N__29782\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31309\,
            in2 => \N__31357\,
            in3 => \N__29770\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__48795\,
            ce => \N__29694\,
            sr => \N__48118\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31332\,
            in2 => \N__31284\,
            in3 => \N__29761\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__48787\,
            ce => \N__29695\,
            sr => \N__48125\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31308\,
            in2 => \N__31260\,
            in3 => \N__29752\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__48787\,
            ce => \N__29695\,
            sr => \N__48125\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31236\,
            in2 => \N__31285\,
            in3 => \N__29743\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__48787\,
            ce => \N__29695\,
            sr => \N__48125\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31095\,
            in2 => \N__31261\,
            in3 => \N__29731\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__48787\,
            ce => \N__29695\,
            sr => \N__48125\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29728\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48787\,
            ce => \N__29695\,
            sr => \N__48125\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__33574\,
            in1 => \N__29995\,
            in2 => \N__33306\,
            in3 => \N__30486\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48779\,
            ce => 'H',
            sr => \N__48129\
        );

    \phase_controller_slave.state_4_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__31008\,
            in1 => \N__45714\,
            in2 => \_gnd_net_\,
            in3 => \N__45923\,
            lcout => \phase_controller_slave.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48770\,
            ce => 'H',
            sr => \N__48134\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__29880\,
            in1 => \N__33780\,
            in2 => \_gnd_net_\,
            in3 => \N__29833\,
            lcout => \current_shift_inst.timer_s1.N_191_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T01_er_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29946\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48754\,
            ce => \N__39520\,
            sr => \N__48147\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42568\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__39875\,
            sr => \N__48153\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42535\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__39875\,
            sr => \N__48153\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39849\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48748\,
            ce => \N__39875\,
            sr => \N__48153\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__46154\,
            in1 => \N__46978\,
            in2 => \N__38998\,
            in3 => \N__43879\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48742\,
            ce => 'H',
            sr => \N__48160\
        );

    \phase_controller_inst1.state_1_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__29977\,
            in1 => \N__39673\,
            in2 => \N__29947\,
            in3 => \N__29905\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48742\,
            ce => 'H',
            sr => \N__48160\
        );

    \current_shift_inst.timer_s1.running_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__29881\,
            in1 => \N__33766\,
            in2 => \_gnd_net_\,
            in3 => \N__29832\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48170\
        );

    \phase_controller_inst1.S1_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39597\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48170\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__46155\,
            in1 => \N__46924\,
            in2 => \N__39038\,
            in3 => \N__43878\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48735\,
            ce => 'H',
            sr => \N__48170\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__49124\,
            in1 => \N__47233\,
            in2 => \_gnd_net_\,
            in3 => \N__46238\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48730\,
            ce => \N__46350\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__46531\,
            in1 => \N__48894\,
            in2 => \N__46167\,
            in3 => \N__46447\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48730\,
            ce => \N__46350\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__46239\,
            in1 => \N__49125\,
            in2 => \_gnd_net_\,
            in3 => \N__47122\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48730\,
            ce => \N__46350\,
            sr => \N__48182\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__49115\,
            in1 => \N__47293\,
            in2 => \_gnd_net_\,
            in3 => \N__46250\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48722\,
            ce => \N__46345\,
            sr => \N__48190\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__46087\,
            in1 => \N__46527\,
            in2 => \N__46166\,
            in3 => \N__46446\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48722\,
            ce => \N__46345\,
            sr => \N__48190\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__32897\,
            in1 => \N__32690\,
            in2 => \N__32570\,
            in3 => \N__30124\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48197\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32526\,
            in1 => \N__32898\,
            in2 => \N__32732\,
            in3 => \N__30112\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48197\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5_3_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__30019\,
            in1 => \N__46569\,
            in2 => \N__38798\,
            in3 => \N__30004\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_14_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__46284\,
            in1 => \N__47427\,
            in2 => \N__36821\,
            in3 => \N__43876\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48197\
        );

    \delay_measurement_inst.delay_tr_reg_15_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__43877\,
            in1 => \N__46285\,
            in2 => \N__38883\,
            in3 => \N__47365\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48715\,
            ce => 'H',
            sr => \N__48197\
        );

    \current_shift_inst.un10_control_input_z_i_31_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34894\,
            lcout => \current_shift_inst.z_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVQKU1_5_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__39994\,
            in1 => \N__39931\,
            in2 => \N__33964\,
            in3 => \N__33914\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVQKU1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_RNIC90O_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31846\,
            in2 => \_gnd_net_\,
            in3 => \N__31760\,
            lcout => \current_shift_inst.timer_phase.N_188_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32402\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_12_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32401\,
            in2 => \_gnd_net_\,
            in3 => \N__32348\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30055\,
            in2 => \N__32317\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_24_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33055\,
            in3 => \N__30049\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30145\,
            in2 => \N__33031\,
            in3 => \N__30139\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33006\,
            in2 => \_gnd_net_\,
            in3 => \N__30136\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32985\,
            in2 => \_gnd_net_\,
            in3 => \N__30133\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32961\,
            in2 => \_gnd_net_\,
            in3 => \N__30130\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32940\,
            in2 => \_gnd_net_\,
            in3 => \N__30127\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32044\,
            in2 => \_gnd_net_\,
            in3 => \N__30115\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32008\,
            in2 => \_gnd_net_\,
            in3 => \N__30103\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_12_25_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_12_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32421\,
            in2 => \_gnd_net_\,
            in3 => \N__30100\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32286\,
            in2 => \_gnd_net_\,
            in3 => \N__30097\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32265\,
            in2 => \_gnd_net_\,
            in3 => \N__30211\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32244\,
            in2 => \_gnd_net_\,
            in3 => \N__30208\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32223\,
            in2 => \_gnd_net_\,
            in3 => \N__30205\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_12_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32202\,
            in2 => \_gnd_net_\,
            in3 => \N__30202\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32145\,
            in3 => \N__30190\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_12_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32442\,
            in2 => \_gnd_net_\,
            in3 => \N__30187\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_12_26_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32181\,
            in2 => \_gnd_net_\,
            in3 => \N__30184\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33075\,
            in2 => \_gnd_net_\,
            in3 => \N__30181\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30178\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111000"
        )
    port map (
            in0 => \N__30523\,
            in1 => \N__33628\,
            in2 => \N__33360\,
            in3 => \N__30484\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48834\,
            ce => 'H',
            sr => \N__48091\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__36063\,
            in1 => \N__30485\,
            in2 => \N__33648\,
            in3 => \N__30357\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48834\,
            ce => 'H',
            sr => \N__48091\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31193\,
            in1 => \N__30335\,
            in2 => \_gnd_net_\,
            in3 => \N__30319\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31205\,
            in1 => \N__30314\,
            in2 => \_gnd_net_\,
            in3 => \N__30298\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31194\,
            in1 => \N__30293\,
            in2 => \_gnd_net_\,
            in3 => \N__30274\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31206\,
            in1 => \N__30269\,
            in2 => \_gnd_net_\,
            in3 => \N__30250\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31195\,
            in1 => \N__30247\,
            in2 => \_gnd_net_\,
            in3 => \N__30232\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31207\,
            in1 => \N__30229\,
            in2 => \_gnd_net_\,
            in3 => \N__30214\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31196\,
            in1 => \N__30725\,
            in2 => \_gnd_net_\,
            in3 => \N__30706\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31208\,
            in1 => \N__30701\,
            in2 => \_gnd_net_\,
            in3 => \N__30682\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__48824\,
            ce => \N__31072\,
            sr => \N__48096\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31216\,
            in1 => \N__30677\,
            in2 => \_gnd_net_\,
            in3 => \N__30658\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31200\,
            in1 => \N__30653\,
            in2 => \_gnd_net_\,
            in3 => \N__30634\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31213\,
            in1 => \N__30629\,
            in2 => \_gnd_net_\,
            in3 => \N__30610\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31197\,
            in1 => \N__30605\,
            in2 => \_gnd_net_\,
            in3 => \N__30586\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31214\,
            in1 => \N__30583\,
            in2 => \_gnd_net_\,
            in3 => \N__30568\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31198\,
            in1 => \N__30565\,
            in2 => \_gnd_net_\,
            in3 => \N__30550\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31215\,
            in1 => \N__30545\,
            in2 => \_gnd_net_\,
            in3 => \N__30526\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31199\,
            in1 => \N__30905\,
            in2 => \_gnd_net_\,
            in3 => \N__30886\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__48814\,
            ce => \N__31082\,
            sr => \N__48104\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31201\,
            in1 => \N__30881\,
            in2 => \_gnd_net_\,
            in3 => \N__30862\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31217\,
            in1 => \N__30857\,
            in2 => \_gnd_net_\,
            in3 => \N__30838\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31202\,
            in1 => \N__30833\,
            in2 => \_gnd_net_\,
            in3 => \N__30814\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31218\,
            in1 => \N__30809\,
            in2 => \_gnd_net_\,
            in3 => \N__30790\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31203\,
            in1 => \N__30787\,
            in2 => \_gnd_net_\,
            in3 => \N__30772\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31219\,
            in1 => \N__30769\,
            in2 => \_gnd_net_\,
            in3 => \N__30754\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31204\,
            in1 => \N__30749\,
            in2 => \_gnd_net_\,
            in3 => \N__30730\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31220\,
            in1 => \N__31355\,
            in2 => \_gnd_net_\,
            in3 => \N__31336\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__48807\,
            ce => \N__31083\,
            sr => \N__48110\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31209\,
            in1 => \N__31331\,
            in2 => \_gnd_net_\,
            in3 => \N__31312\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__48796\,
            ce => \N__31084\,
            sr => \N__48119\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31221\,
            in1 => \N__31307\,
            in2 => \_gnd_net_\,
            in3 => \N__31288\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__48796\,
            ce => \N__31084\,
            sr => \N__48119\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31210\,
            in1 => \N__31283\,
            in2 => \_gnd_net_\,
            in3 => \N__31264\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__48796\,
            ce => \N__31084\,
            sr => \N__48119\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31222\,
            in1 => \N__31259\,
            in2 => \_gnd_net_\,
            in3 => \N__31240\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__48796\,
            ce => \N__31084\,
            sr => \N__48119\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31211\,
            in1 => \N__31237\,
            in2 => \_gnd_net_\,
            in3 => \N__31225\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__48796\,
            ce => \N__31084\,
            sr => \N__48119\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31096\,
            in1 => \N__31212\,
            in2 => \_gnd_net_\,
            in3 => \N__31099\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48796\,
            ce => \N__31084\,
            sr => \N__48119\
        );

    \phase_controller_slave.state_RNO_0_3_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__30992\,
            in1 => \N__45713\,
            in2 => \_gnd_net_\,
            in3 => \N__45922\,
            lcout => \phase_controller_slave.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39853\,
            lcout => \current_shift_inst.elapsed_time_ns_1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48772\,
            ce => \N__39878\,
            sr => \N__48135\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__42230\,
            in1 => \N__41978\,
            in2 => \N__42196\,
            in3 => \N__42600\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__31464\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__42601\,
            in1 => \N__42191\,
            in2 => \N__42002\,
            in3 => \N__42231\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__31464\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__45433\,
            in1 => \N__45361\,
            in2 => \N__45655\,
            in3 => \N__45872\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__31464\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__45873\,
            in1 => \N__45643\,
            in2 => \N__45391\,
            in3 => \N__45434\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__31464\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__43987\,
            in1 => \N__44006\,
            in2 => \_gnd_net_\,
            in3 => \N__43951\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48762\,
            ce => \N__31464\,
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31387\,
            lcout => \current_shift_inst.un4_control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31381\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38743\,
            lcout => \current_shift_inst.un4_control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIN7DV_8_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40632\,
            in2 => \_gnd_net_\,
            in3 => \N__34468\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIN7DV_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4H5J_19_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40911\,
            in2 => \_gnd_net_\,
            in3 => \N__34708\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4H5J_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDLO51_11_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__34339\,
            in1 => \N__40340\,
            in2 => \N__40423\,
            in3 => \N__34303\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDLO51_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIU73K_23_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41662\,
            in2 => \_gnd_net_\,
            in3 => \N__34549\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIU73K_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIJTQ51_12_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__40269\,
            in1 => \N__40341\,
            in2 => \N__34311\,
            in3 => \N__34258\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJTQ51_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIVDV51_14_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40193\,
            in1 => \N__34861\,
            in2 => \N__34233\,
            in3 => \N__41183\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIVDV51_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIPC571_19_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__40912\,
            in1 => \N__40838\,
            in2 => \N__34718\,
            in3 => \N__34669\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPC571_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBU361_16_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__34819\,
            in1 => \N__41043\,
            in2 => \N__41116\,
            in3 => \N__34784\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBU361_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_RNO_0_25_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110010110"
        )
    port map (
            in0 => \N__41890\,
            in1 => \N__37408\,
            in2 => \N__41851\,
            in3 => \N__34913\,
            lcout => \current_shift_inst.un38_control_input_0_axb_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI4D1J_16_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41115\,
            in2 => \_gnd_net_\,
            in3 => \N__34833\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI4D1J_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIHCE81_26_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__41469\,
            in1 => \N__41405\,
            in2 => \N__35056\,
            in3 => \N__35024\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIHCE81_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.running_RNIL91O_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__31791\,
            in1 => \N__31845\,
            in2 => \_gnd_net_\,
            in3 => \N__31761\,
            lcout => \current_shift_inst.timer_phase.N_192_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7K6K_26_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41468\,
            in2 => \_gnd_net_\,
            in3 => \N__35050\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7K6K_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIAO7K_27_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41406\,
            in2 => \_gnd_net_\,
            in3 => \N__35023\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIAO7K_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIDS8K_28_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41338\,
            in2 => \_gnd_net_\,
            in3 => \N__34985\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIDS8K_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_RNIMR6L_0_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__43947\,
            in1 => \N__43981\,
            in2 => \_gnd_net_\,
            in3 => \N__44010\,
            lcout => \delay_measurement_inst.tr_state_RNIMR6LZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5S981_24_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__35117\,
            in1 => \N__41526\,
            in2 => \N__41590\,
            in3 => \N__35080\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5S981_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIB4C81_25_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__41527\,
            in1 => \N__41470\,
            in2 => \N__35090\,
            in3 => \N__35054\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIB4C81_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNINKG81_27_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__41407\,
            in1 => \N__41337\,
            in2 => \N__35029\,
            in3 => \N__34984\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINKG81_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNIBBPU1_7_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__34515\,
            in1 => \N__40628\,
            in2 => \N__40705\,
            in3 => \N__34479\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIBBPU1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__46382\,
            in1 => \N__39164\,
            in2 => \N__39122\,
            in3 => \N__39080\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48731\,
            ce => \N__46641\,
            sr => \N__48183\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__39286\,
            in1 => \N__39165\,
            in2 => \N__39261\,
            in3 => \N__39079\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48731\,
            ce => \N__46641\,
            sr => \N__48183\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__39081\,
            in1 => \N__39112\,
            in2 => \_gnd_net_\,
            in3 => \N__39166\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48731\,
            ce => \N__46641\,
            sr => \N__48183\
        );

    \current_shift_inst.timer_phase.running_RNIB31B_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31844\,
            lcout => \current_shift_inst.timer_phase.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__45134\,
            in1 => \N__45053\,
            in2 => \N__38799\,
            in3 => \N__45006\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000001"
        )
    port map (
            in0 => \N__45007\,
            in1 => \N__45135\,
            in2 => \N__45058\,
            in3 => \N__38962\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__45136\,
            in1 => \N__39003\,
            in2 => \_gnd_net_\,
            in3 => \N__45004\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39832\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__39037\,
            in1 => \N__45133\,
            in2 => \_gnd_net_\,
            in3 => \N__45005\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__45132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38869\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__38867\,
            in1 => \N__45131\,
            in2 => \_gnd_net_\,
            in3 => \N__36811\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__36973\,
            in1 => \N__38868\,
            in2 => \N__39220\,
            in3 => \N__38833\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48724\,
            ce => \N__46628\,
            sr => \N__48191\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31927\,
            in2 => \N__31942\,
            in3 => \N__32316\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_13_21_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31909\,
            in2 => \N__31921\,
            in3 => \N__33054\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31891\,
            in2 => \N__31903\,
            in3 => \N__33030\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31885\,
            in2 => \N__46666\,
            in3 => \N__33007\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31870\,
            in2 => \N__31879\,
            in3 => \N__32986\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31852\,
            in2 => \N__31864\,
            in3 => \N__32965\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32941\,
            in1 => \N__32059\,
            in2 => \N__32068\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32026\,
            in2 => \N__32053\,
            in3 => \N__32043\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31990\,
            in2 => \N__32020\,
            in3 => \N__32007\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31984\,
            in2 => \N__37057\,
            in3 => \N__32422\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31978\,
            in2 => \N__37042\,
            in3 => \N__32287\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31972\,
            in2 => \N__37027\,
            in3 => \N__32266\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31966\,
            in2 => \N__36952\,
            in3 => \N__32245\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31948\,
            in2 => \N__31960\,
            in3 => \N__32224\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32152\,
            in2 => \N__32167\,
            in3 => \N__32203\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32125\,
            in2 => \N__44035\,
            in3 => \N__32146\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32119\,
            in2 => \N__32086\,
            in3 => \N__32443\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32101\,
            in2 => \N__32113\,
            in3 => \N__32182\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32095\,
            in2 => \N__32077\,
            in3 => \N__33076\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32089\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39786\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48708\,
            ce => \N__46642\,
            sr => \N__48211\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39740\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48708\,
            ce => \N__46642\,
            sr => \N__48211\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32899\,
            in1 => \N__32573\,
            in2 => \N__32777\,
            in3 => \N__32428\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__32407\,
            in1 => \N__32315\,
            in2 => \_gnd_net_\,
            in3 => \N__32350\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000011010000"
        )
    port map (
            in0 => \N__32902\,
            in1 => \N__32576\,
            in2 => \N__32320\,
            in3 => \N__32757\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__32293\,
            in1 => \N__32758\,
            in2 => \N__32594\,
            in3 => \N__32903\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32900\,
            in1 => \N__32574\,
            in2 => \N__32778\,
            in3 => \N__32272\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32571\,
            in1 => \N__32759\,
            in2 => \N__32925\,
            in3 => \N__32251\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32901\,
            in1 => \N__32575\,
            in2 => \N__32779\,
            in3 => \N__32230\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32572\,
            in1 => \N__32760\,
            in2 => \N__32926\,
            in3 => \N__32209\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48705\,
            ce => 'H',
            sr => \N__48216\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32581\,
            in1 => \N__32907\,
            in2 => \N__32773\,
            in3 => \N__32188\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32904\,
            in1 => \N__32584\,
            in2 => \N__32770\,
            in3 => \N__33082\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010100010"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__32737\,
            in2 => \N__32595\,
            in3 => \N__32913\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_13_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010000010"
        )
    port map (
            in0 => \N__33037\,
            in1 => \N__32744\,
            in2 => \N__32923\,
            in3 => \N__32590\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_13_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32582\,
            in1 => \N__32908\,
            in2 => \N__32774\,
            in3 => \N__33013\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_13_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32905\,
            in1 => \N__32585\,
            in2 => \N__32771\,
            in3 => \N__32992\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__32583\,
            in1 => \N__32909\,
            in2 => \N__32775\,
            in3 => \N__32971\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__32906\,
            in1 => \N__32586\,
            in2 => \N__32772\,
            in3 => \N__32947\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48703\,
            ce => 'H',
            sr => \N__48222\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_13_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__32924\,
            in1 => \N__32785\,
            in2 => \N__32776\,
            in3 => \N__32580\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48701\,
            ce => 'H',
            sr => \N__48224\
        );

    \phase_controller_inst1.S2_LC_13_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39694\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48700\,
            ce => 'H',
            sr => \N__48229\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__42270\,
            in1 => \N__42042\,
            in2 => \N__42195\,
            in3 => \N__44845\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48825\,
            ce => 'H',
            sr => \N__48097\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__33632\,
            in1 => \N__36339\,
            in2 => \_gnd_net_\,
            in3 => \N__33455\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48825\,
            ce => 'H',
            sr => \N__48097\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36319\,
            in1 => \N__33412\,
            in2 => \_gnd_net_\,
            in3 => \N__36646\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48815\,
            ce => \N__36226\,
            sr => \N__48105\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__36584\,
            in1 => \_gnd_net_\,
            in2 => \N__36367\,
            in3 => \N__33364\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48808\,
            ce => \N__36231\,
            sr => \N__48111\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__33309\,
            in1 => \N__36344\,
            in2 => \_gnd_net_\,
            in3 => \N__36585\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48808\,
            ce => \N__36231\,
            sr => \N__48111\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__36586\,
            in1 => \_gnd_net_\,
            in2 => \N__36368\,
            in3 => \N__33259\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48808\,
            ce => \N__36231\,
            sr => \N__48111\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__33211\,
            in1 => \N__36348\,
            in2 => \_gnd_net_\,
            in3 => \N__36587\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48808\,
            ce => \N__36231\,
            sr => \N__48111\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__36340\,
            in1 => \N__33163\,
            in2 => \_gnd_net_\,
            in3 => \N__33129\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48808\,
            ce => \N__36231\,
            sr => \N__48111\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45456\,
            in2 => \_gnd_net_\,
            in3 => \N__45365\,
            lcout => \phase_controller_slave.stoper_tr.time_passed11\,
            ltout => \phase_controller_slave.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33691\,
            in3 => \N__45870\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33688\,
            in2 => \N__38407\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38380\,
            in2 => \_gnd_net_\,
            in3 => \N__33682\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33790\,
            in2 => \N__38362\,
            in3 => \N__33679\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38329\,
            in2 => \_gnd_net_\,
            in3 => \N__33676\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38311\,
            in2 => \_gnd_net_\,
            in3 => \N__33673\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38281\,
            in2 => \_gnd_net_\,
            in3 => \N__33670\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38251\,
            in2 => \_gnd_net_\,
            in3 => \N__33667\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38218\,
            in2 => \_gnd_net_\,
            in3 => \N__33718\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38611\,
            in2 => \_gnd_net_\,
            in3 => \N__33715\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38581\,
            in3 => \N__33712\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45778\,
            in2 => \_gnd_net_\,
            in3 => \N__33709\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38524\,
            in2 => \_gnd_net_\,
            in3 => \N__33706\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38506\,
            in3 => \N__33703\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38458\,
            in2 => \_gnd_net_\,
            in3 => \N__33700\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38425\,
            in2 => \_gnd_net_\,
            in3 => \N__33697\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38734\,
            in2 => \_gnd_net_\,
            in3 => \N__33694\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38713\,
            in2 => \_gnd_net_\,
            in3 => \N__33799\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38695\,
            in3 => \N__33796\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38674\,
            in2 => \_gnd_net_\,
            in3 => \N__33793\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45900\,
            in2 => \_gnd_net_\,
            in3 => \N__45861\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42219\,
            in2 => \_gnd_net_\,
            in3 => \N__41967\,
            lcout => \phase_controller_slave.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33779\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_RNI48NB_31_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33742\,
            in2 => \N__34143\,
            in3 => \N__34136\,
            lcout => \current_shift_inst.un38_control_input_0\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_1_c_RNIJF2G_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33736\,
            in2 => \_gnd_net_\,
            in3 => \N__33730\,
            lcout => \current_shift_inst.un4_control_input_cry_1_c_RNIJF2GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_1\,
            carryout => \current_shift_inst.un4_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_2_c_RNILI3G_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33727\,
            in2 => \_gnd_net_\,
            in3 => \N__33721\,
            lcout => \current_shift_inst.un4_control_input_cry_2_c_RNILI3GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_2\,
            carryout => \current_shift_inst.un4_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_3_c_RNINL4G_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36784\,
            in2 => \_gnd_net_\,
            in3 => \N__33826\,
            lcout => \current_shift_inst.un4_control_input_cry_3_c_RNINL4GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_3\,
            carryout => \current_shift_inst.un4_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_4_c_RNIPO5G_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36778\,
            in2 => \_gnd_net_\,
            in3 => \N__33823\,
            lcout => \current_shift_inst.un4_control_input_cry_4_c_RNIPO5GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_4\,
            carryout => \current_shift_inst.un4_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_5_c_RNIRR6G_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36874\,
            in2 => \_gnd_net_\,
            in3 => \N__33820\,
            lcout => \current_shift_inst.un4_control_input_cry_5_c_RNIRR6GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_5\,
            carryout => \current_shift_inst.un4_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_6_c_RNITU7G_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36868\,
            in2 => \_gnd_net_\,
            in3 => \N__33817\,
            lcout => \current_shift_inst.un4_control_input_cry_6_c_RNITU7GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_6\,
            carryout => \current_shift_inst.un4_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_7_c_RNIV19G_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36862\,
            in2 => \_gnd_net_\,
            in3 => \N__33814\,
            lcout => \current_shift_inst.un4_control_input_cry_7_c_RNIV19GZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_7\,
            carryout => \current_shift_inst.un4_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_8_c_RNI15AG_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36856\,
            in2 => \_gnd_net_\,
            in3 => \N__33811\,
            lcout => \current_shift_inst.un4_control_input_cry_8_c_RNI15AGZ0\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_9_c_RNIALDJ_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36850\,
            in2 => \_gnd_net_\,
            in3 => \N__33808\,
            lcout => \current_shift_inst.un4_control_input_cry_9_c_RNIALDJZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_9\,
            carryout => \current_shift_inst.un4_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_10_c_RNIJLTG_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36844\,
            in2 => \_gnd_net_\,
            in3 => \N__33805\,
            lcout => \current_shift_inst.un4_control_input_cry_10_c_RNIJLTGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_10\,
            carryout => \current_shift_inst.un4_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_11_c_RNILOUG_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36934\,
            in2 => \_gnd_net_\,
            in3 => \N__33802\,
            lcout => \current_shift_inst.un4_control_input_cry_11_c_RNILOUGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_11\,
            carryout => \current_shift_inst.un4_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_12_c_RNINRVG_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37192\,
            in2 => \_gnd_net_\,
            in3 => \N__33853\,
            lcout => \current_shift_inst.un4_control_input_cry_12_c_RNINRVGZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_12\,
            carryout => \current_shift_inst.un4_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_13_c_RNIPU0H_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43525\,
            in2 => \_gnd_net_\,
            in3 => \N__33850\,
            lcout => \current_shift_inst.un4_control_input_cry_13_c_RNIPU0HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_13\,
            carryout => \current_shift_inst.un4_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_14_c_RNIR12H_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36916\,
            in3 => \N__33847\,
            lcout => \current_shift_inst.un4_control_input_cry_14_c_RNIR12HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_14\,
            carryout => \current_shift_inst.un4_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_15_c_RNIT43H_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36907\,
            in3 => \N__33844\,
            lcout => \current_shift_inst.un4_control_input_cry_15_c_RNIT43HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_15\,
            carryout => \current_shift_inst.un4_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_16_c_RNIV74H_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36922\,
            in2 => \_gnd_net_\,
            in3 => \N__33841\,
            lcout => \current_shift_inst.un4_control_input_cry_16_c_RNIV74HZ0\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_17_c_RNI1B5H_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36898\,
            in2 => \_gnd_net_\,
            in3 => \N__33838\,
            lcout => \current_shift_inst.un4_control_input_cry_17_c_RNI1B5HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_17\,
            carryout => \current_shift_inst.un4_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_18_c_RNI3E6H_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36928\,
            in2 => \_gnd_net_\,
            in3 => \N__33835\,
            lcout => \current_shift_inst.un4_control_input_cry_18_c_RNI3E6HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_18\,
            carryout => \current_shift_inst.un4_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_19_c_RNIS88H_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36880\,
            in2 => \_gnd_net_\,
            in3 => \N__33832\,
            lcout => \current_shift_inst.un4_control_input_cry_19_c_RNIS88HZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_19\,
            carryout => \current_shift_inst.un4_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_20_c_RNILQ1I_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37201\,
            in2 => \_gnd_net_\,
            in3 => \N__33829\,
            lcout => \current_shift_inst.un4_control_input_cry_20_c_RNILQ1IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_20\,
            carryout => \current_shift_inst.un4_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_21_c_RNINT2I_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36838\,
            in2 => \_gnd_net_\,
            in3 => \N__33880\,
            lcout => \current_shift_inst.un4_control_input_cry_21_c_RNINT2IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_21\,
            carryout => \current_shift_inst.un4_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_22_c_RNIP04I_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36892\,
            in2 => \_gnd_net_\,
            in3 => \N__33877\,
            lcout => \current_shift_inst.un4_control_input_cry_22_c_RNIP04IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_22\,
            carryout => \current_shift_inst.un4_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_23_c_RNIR35I_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43510\,
            in2 => \_gnd_net_\,
            in3 => \N__33874\,
            lcout => \current_shift_inst.un4_control_input_cry_23_c_RNIR35IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_23\,
            carryout => \current_shift_inst.un4_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_24_c_RNIT66I_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37063\,
            in2 => \_gnd_net_\,
            in3 => \N__33871\,
            lcout => \current_shift_inst.un4_control_input_cry_24_c_RNIT66IZ0\,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.un4_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_25_c_RNIV97I_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37081\,
            in2 => \_gnd_net_\,
            in3 => \N__33868\,
            lcout => \current_shift_inst.un4_control_input_cry_25_c_RNIV97IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_25\,
            carryout => \current_shift_inst.un4_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_26_c_RNI1D8I_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36886\,
            in2 => \_gnd_net_\,
            in3 => \N__33865\,
            lcout => \current_shift_inst.un4_control_input_cry_26_c_RNI1D8IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_26\,
            carryout => \current_shift_inst.un4_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_27_c_RNI3G9I_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37069\,
            in2 => \_gnd_net_\,
            in3 => \N__33862\,
            lcout => \current_shift_inst.un4_control_input_cry_27_c_RNI3G9IZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_27\,
            carryout => \current_shift_inst.un4_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_28_c_RNI5JAI_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37075\,
            in2 => \_gnd_net_\,
            in3 => \N__33859\,
            lcout => \current_shift_inst.un4_control_input_cry_28_c_RNI5JAIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_28\,
            carryout => \current_shift_inst.un4_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_29_c_RNIUDCI_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37087\,
            in2 => \_gnd_net_\,
            in3 => \N__33856\,
            lcout => \current_shift_inst.un4_control_input_cry_29_c_RNIUDCIZ0\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_cry_29\,
            carryout => \current_shift_inst.un4_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_cry_30_c_RNINV5J_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37409\,
            in2 => \_gnd_net_\,
            in3 => \N__34192\,
            lcout => \current_shift_inst.un4_control_input_cry_30_c_RNINV5JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI7H2J_17_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41036\,
            in2 => \_gnd_net_\,
            in3 => \N__34783\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI7H2J_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_0_c_inv_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34161\,
            in2 => \N__34117\,
            in3 => \N__34144\,
            lcout => \G_407\,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.z_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_1_c_inv_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34095\,
            in2 => \N__34078\,
            in3 => \N__37328\,
            lcout => \G_406\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_0\,
            carryout => \current_shift_inst.z_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_2_c_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37267\,
            in2 => \N__34058\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_1\,
            carryout => \current_shift_inst.z_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_3_c_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37255\,
            in2 => \N__34032\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_2\,
            carryout => \current_shift_inst.z_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_4_c_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33989\,
            in2 => \N__37243\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_3\,
            carryout => \current_shift_inst.z_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_5_c_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37228\,
            in2 => \N__33943\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_4\,
            carryout => \current_shift_inst.z_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_6_c_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33897\,
            in2 => \N__37216\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_5\,
            carryout => \current_shift_inst.z_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_7_c_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34505\,
            in2 => \N__37582\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_6\,
            carryout => \current_shift_inst.z_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_8_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37564\,
            in2 => \N__34478\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.z_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_9_c_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34421\,
            in2 => \N__37549\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_8\,
            carryout => \current_shift_inst.z_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_10_c_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37534\,
            in2 => \N__34393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_9\,
            carryout => \current_shift_inst.z_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_11_c_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37522\,
            in2 => \N__34356\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_10\,
            carryout => \current_shift_inst.z_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_12_c_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34307\,
            in2 => \N__37510\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_11\,
            carryout => \current_shift_inst.z_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_13_c_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37495\,
            in2 => \N__34268\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_12\,
            carryout => \current_shift_inst.z_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_14_c_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34219\,
            in2 => \N__37483\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_13\,
            carryout => \current_shift_inst.z_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_15_c_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34865\,
            in2 => \N__37705\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_14\,
            carryout => \current_shift_inst.z_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_16_c_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34829\,
            in2 => \N__37687\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.z_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_17_c_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37669\,
            in2 => \N__34794\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_16\,
            carryout => \current_shift_inst.z_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_18_c_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34748\,
            in2 => \N__37654\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_17\,
            carryout => \current_shift_inst.z_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_19_c_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37636\,
            in2 => \N__34722\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_18\,
            carryout => \current_shift_inst.z_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_20_c_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37624\,
            in2 => \N__34687\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_19\,
            carryout => \current_shift_inst.z_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_21_c_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37609\,
            in2 => \N__34635\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_20\,
            carryout => \current_shift_inst.z_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_22_c_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37597\,
            in2 => \N__34594\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_21\,
            carryout => \current_shift_inst.z_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_23_c_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34550\,
            in2 => \N__37855\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_22\,
            carryout => \current_shift_inst.z_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_24_c_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35118\,
            in2 => \N__37837\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_21_0_\,
            carryout => \current_shift_inst.z_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_25_c_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37819\,
            in2 => \N__35091\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_24\,
            carryout => \current_shift_inst.z_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_26_c_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35055\,
            in2 => \N__37804\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_25\,
            carryout => \current_shift_inst.z_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_27_c_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35028\,
            in2 => \N__37786\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_26\,
            carryout => \current_shift_inst.z_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_28_c_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37768\,
            in2 => \N__35001\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_27\,
            carryout => \current_shift_inst.z_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_29_c_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34958\,
            in2 => \N__37753\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_28\,
            carryout => \current_shift_inst.z_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_cry_30_c_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37735\,
            in2 => \N__34926\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.z_cry_29\,
            carryout => \current_shift_inst.z_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_s_31_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__37427\,
            in1 => \N__37717\,
            in2 => \N__41847\,
            in3 => \N__34897\,
            lcout => \current_shift_inst.z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.counter_0_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35584\,
            in1 => \N__40118\,
            in2 => \_gnd_net_\,
            in3 => \N__35158\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_22_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_0\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_1_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35579\,
            in1 => \N__40083\,
            in2 => \_gnd_net_\,
            in3 => \N__35155\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_0\,
            carryout => \current_shift_inst.timer_phase.counter_cry_1\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_2_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35585\,
            in1 => \N__40016\,
            in2 => \_gnd_net_\,
            in3 => \N__35152\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_1\,
            carryout => \current_shift_inst.timer_phase.counter_cry_2\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_3_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35580\,
            in1 => \N__39953\,
            in2 => \_gnd_net_\,
            in3 => \N__35149\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_2\,
            carryout => \current_shift_inst.timer_phase.counter_cry_3\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_4_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35586\,
            in1 => \N__40721\,
            in2 => \_gnd_net_\,
            in3 => \N__35146\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_3\,
            carryout => \current_shift_inst.timer_phase.counter_cry_4\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_5_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35581\,
            in1 => \N__40652\,
            in2 => \_gnd_net_\,
            in3 => \N__35143\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_4\,
            carryout => \current_shift_inst.timer_phase.counter_cry_5\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_6_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35583\,
            in1 => \N__40580\,
            in2 => \_gnd_net_\,
            in3 => \N__35140\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_5\,
            carryout => \current_shift_inst.timer_phase.counter_cry_6\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_7_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35582\,
            in1 => \N__40520\,
            in2 => \_gnd_net_\,
            in3 => \N__35137\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_6\,
            carryout => \current_shift_inst.timer_phase.counter_cry_7\,
            clk => \N__48717\,
            ce => \N__35480\,
            sr => \N__48198\
        );

    \current_shift_inst.timer_phase.counter_8_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35590\,
            in1 => \N__40442\,
            in2 => \_gnd_net_\,
            in3 => \N__35134\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_23_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_8\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_9_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35594\,
            in1 => \N__40358\,
            in2 => \_gnd_net_\,
            in3 => \N__35185\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_8\,
            carryout => \current_shift_inst.timer_phase.counter_cry_9\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_10_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35587\,
            in1 => \N__40298\,
            in2 => \_gnd_net_\,
            in3 => \N__35182\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_9\,
            carryout => \current_shift_inst.timer_phase.counter_cry_10\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_11_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35591\,
            in1 => \N__40217\,
            in2 => \_gnd_net_\,
            in3 => \N__35179\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_10\,
            carryout => \current_shift_inst.timer_phase.counter_cry_11\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_12_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35588\,
            in1 => \N__41207\,
            in2 => \_gnd_net_\,
            in3 => \N__35176\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_11\,
            carryout => \current_shift_inst.timer_phase.counter_cry_12\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_13_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35592\,
            in1 => \N__41132\,
            in2 => \_gnd_net_\,
            in3 => \N__35173\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_12\,
            carryout => \current_shift_inst.timer_phase.counter_cry_13\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_14_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35589\,
            in1 => \N__41063\,
            in2 => \_gnd_net_\,
            in3 => \N__35170\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_13\,
            carryout => \current_shift_inst.timer_phase.counter_cry_14\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_15_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35593\,
            in1 => \N__41000\,
            in2 => \_gnd_net_\,
            in3 => \N__35167\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_14\,
            carryout => \current_shift_inst.timer_phase.counter_cry_15\,
            clk => \N__48711\,
            ce => \N__35476\,
            sr => \N__48206\
        );

    \current_shift_inst.timer_phase.counter_16_LC_14_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35595\,
            in1 => \N__40928\,
            in2 => \_gnd_net_\,
            in3 => \N__35164\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_24_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_16\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_17_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35601\,
            in1 => \N__40862\,
            in2 => \_gnd_net_\,
            in3 => \N__35161\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_16\,
            carryout => \current_shift_inst.timer_phase.counter_cry_17\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_18_LC_14_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35596\,
            in1 => \N__40793\,
            in2 => \_gnd_net_\,
            in3 => \N__35212\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_17\,
            carryout => \current_shift_inst.timer_phase.counter_cry_18\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_19_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35602\,
            in1 => \N__41750\,
            in2 => \_gnd_net_\,
            in3 => \N__35209\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_18\,
            carryout => \current_shift_inst.timer_phase.counter_cry_19\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_20_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35597\,
            in1 => \N__41678\,
            in2 => \_gnd_net_\,
            in3 => \N__35206\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_19\,
            carryout => \current_shift_inst.timer_phase.counter_cry_20\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_21_LC_14_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35603\,
            in1 => \N__41606\,
            in2 => \_gnd_net_\,
            in3 => \N__35203\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_20\,
            carryout => \current_shift_inst.timer_phase.counter_cry_21\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_22_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35598\,
            in1 => \N__41546\,
            in2 => \_gnd_net_\,
            in3 => \N__35200\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_21\,
            carryout => \current_shift_inst.timer_phase.counter_cry_22\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_23_LC_14_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35604\,
            in1 => \N__41484\,
            in2 => \_gnd_net_\,
            in3 => \N__35197\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_22\,
            carryout => \current_shift_inst.timer_phase.counter_cry_23\,
            clk => \N__48709\,
            ce => \N__35481\,
            sr => \N__48212\
        );

    \current_shift_inst.timer_phase.counter_24_LC_14_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35605\,
            in1 => \N__41426\,
            in2 => \_gnd_net_\,
            in3 => \N__35194\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_25_0_\,
            carryout => \current_shift_inst.timer_phase.counter_cry_24\,
            clk => \N__48706\,
            ce => \N__35482\,
            sr => \N__48217\
        );

    \current_shift_inst.timer_phase.counter_25_LC_14_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35599\,
            in1 => \N__41354\,
            in2 => \_gnd_net_\,
            in3 => \N__35191\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_24\,
            carryout => \current_shift_inst.timer_phase.counter_cry_25\,
            clk => \N__48706\,
            ce => \N__35482\,
            sr => \N__48217\
        );

    \current_shift_inst.timer_phase.counter_26_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35606\,
            in1 => \N__41270\,
            in2 => \_gnd_net_\,
            in3 => \N__35188\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_25\,
            carryout => \current_shift_inst.timer_phase.counter_cry_26\,
            clk => \N__48706\,
            ce => \N__35482\,
            sr => \N__48217\
        );

    \current_shift_inst.timer_phase.counter_27_LC_14_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35600\,
            in1 => \N__41927\,
            in2 => \_gnd_net_\,
            in3 => \N__35614\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_26\,
            carryout => \current_shift_inst.timer_phase.counter_cry_27\,
            clk => \N__48706\,
            ce => \N__35482\,
            sr => \N__48217\
        );

    \current_shift_inst.timer_phase.counter_28_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__41286\,
            in2 => \_gnd_net_\,
            in3 => \N__35611\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.counter_cry_27\,
            carryout => \current_shift_inst.timer_phase.counter_cry_28\,
            clk => \N__48706\,
            ce => \N__35482\,
            sr => \N__48217\
        );

    \current_shift_inst.timer_phase.counter_29_LC_14_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__41904\,
            in1 => \N__35608\,
            in2 => \_gnd_net_\,
            in3 => \N__35485\,
            lcout => \current_shift_inst.timer_phase.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48706\,
            ce => \N__35482\,
            sr => \N__48217\
        );

    \SB_DFF_inst_DELAY_TR1_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35443\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR2_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35434\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36667\,
            in1 => \N__36335\,
            in2 => \_gnd_net_\,
            in3 => \N__35428\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48840\,
            ce => \N__36222\,
            sr => \N__48089\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__36663\,
            in1 => \N__36315\,
            in2 => \N__35801\,
            in3 => \N__35374\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48835\,
            ce => \N__36232\,
            sr => \N__48092\
        );

    \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__35319\,
            in1 => \N__35791\,
            in2 => \N__36357\,
            in3 => \N__36661\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48835\,
            ce => \N__36232\,
            sr => \N__48092\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__36665\,
            in1 => \N__36317\,
            in2 => \N__35803\,
            in3 => \N__35265\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48835\,
            ce => \N__36232\,
            sr => \N__48092\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36318\,
            in1 => \N__36151\,
            in2 => \_gnd_net_\,
            in3 => \N__36666\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48835\,
            ce => \N__36232\,
            sr => \N__48092\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__36664\,
            in1 => \N__36316\,
            in2 => \N__35802\,
            in3 => \N__36085\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48835\,
            ce => \N__36232\,
            sr => \N__48092\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__36314\,
            in1 => \N__36031\,
            in2 => \_gnd_net_\,
            in3 => \N__36662\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48835\,
            ce => \N__36232\,
            sr => \N__48092\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__36653\,
            in1 => \N__35983\,
            in2 => \N__36361\,
            in3 => \N__35780\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35932\,
            in1 => \N__36321\,
            in2 => \_gnd_net_\,
            in3 => \N__36648\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__36649\,
            in1 => \_gnd_net_\,
            in2 => \N__36358\,
            in3 => \N__35890\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.target_time_0_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35778\,
            in1 => \N__36320\,
            in2 => \N__35848\,
            in3 => \N__36647\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__36651\,
            in1 => \N__35779\,
            in2 => \N__36359\,
            in3 => \N__35708\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35668\,
            in1 => \N__36325\,
            in2 => \_gnd_net_\,
            in3 => \N__36650\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000001000"
        )
    port map (
            in0 => \N__36652\,
            in1 => \N__36491\,
            in2 => \N__36360\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48826\,
            ce => \N__36227\,
            sr => \N__48098\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42005\,
            in1 => \N__42152\,
            in2 => \N__42306\,
            in3 => \N__44227\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48816\,
            ce => 'H',
            sr => \N__48106\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42006\,
            in1 => \N__42153\,
            in2 => \N__42307\,
            in3 => \N__44710\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48816\,
            ce => 'H',
            sr => \N__48106\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__42151\,
            in1 => \_gnd_net_\,
            in2 => \N__42271\,
            in3 => \N__42004\,
            lcout => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__45896\,
            in1 => \N__38406\,
            in2 => \_gnd_net_\,
            in3 => \N__45871\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__45626\,
            in1 => \N__45458\,
            in2 => \N__36235\,
            in3 => \N__45374\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48816\,
            ce => 'H',
            sr => \N__48106\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__42003\,
            in1 => \N__42150\,
            in2 => \_gnd_net_\,
            in3 => \N__42250\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__45625\,
            in1 => \N__45457\,
            in2 => \N__45394\,
            in3 => \N__36178\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48816\,
            ce => 'H',
            sr => \N__48106\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45507\,
            in1 => \N__45390\,
            in2 => \N__45650\,
            in3 => \N__36169\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45384\,
            in1 => \N__45512\,
            in2 => \N__36160\,
            in3 => \N__45619\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__45508\,
            in1 => \N__36736\,
            in2 => \N__45647\,
            in3 => \N__45387\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45385\,
            in1 => \N__45513\,
            in2 => \N__36730\,
            in3 => \N__45620\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__45509\,
            in1 => \N__36721\,
            in2 => \N__45648\,
            in3 => \N__45388\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45386\,
            in1 => \N__45514\,
            in2 => \N__36715\,
            in3 => \N__45621\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010000100"
        )
    port map (
            in0 => \N__45510\,
            in1 => \N__36706\,
            in2 => \N__45649\,
            in3 => \N__45389\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45383\,
            in1 => \N__45511\,
            in2 => \N__36700\,
            in3 => \N__45618\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48809\,
            ce => 'H',
            sr => \N__48112\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45378\,
            in1 => \N__45630\,
            in2 => \N__36691\,
            in3 => \N__45506\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45499\,
            in1 => \N__45379\,
            in2 => \N__45651\,
            in3 => \N__36682\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45375\,
            in1 => \N__45627\,
            in2 => \N__36676\,
            in3 => \N__45503\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45500\,
            in1 => \N__45380\,
            in2 => \N__45652\,
            in3 => \N__36772\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45376\,
            in1 => \N__45628\,
            in2 => \N__36766\,
            in3 => \N__45504\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45501\,
            in1 => \N__45381\,
            in2 => \N__45653\,
            in3 => \N__36757\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__45377\,
            in1 => \N__45629\,
            in2 => \N__36751\,
            in3 => \N__45505\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__45502\,
            in1 => \N__45382\,
            in2 => \N__45654\,
            in3 => \N__36742\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48797\,
            ce => 'H',
            sr => \N__48120\
        );

    \phase_controller_slave.stoper_tr.target_time_6_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000101"
        )
    port map (
            in0 => \N__45034\,
            in1 => \N__38955\,
            in2 => \N__45165\,
            in3 => \N__44974\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__45212\,
            sr => \N__48126\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__44973\,
            in1 => \N__45157\,
            in2 => \N__46570\,
            in3 => \N__45033\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__45212\,
            sr => \N__48126\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__39004\,
            in1 => \_gnd_net_\,
            in2 => \N__45166\,
            in3 => \N__44972\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__45212\,
            sr => \N__48126\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100010001"
        )
    port map (
            in0 => \N__38896\,
            in1 => \N__36828\,
            in2 => \N__39219\,
            in3 => \N__38825\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__45164\,
            in1 => \_gnd_net_\,
            in2 => \N__36832\,
            in3 => \N__39045\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__45212\,
            sr => \N__48126\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110001"
        )
    port map (
            in0 => \N__38826\,
            in1 => \N__37011\,
            in2 => \N__38912\,
            in3 => \N__39214\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__45212\,
            sr => \N__48126\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__38897\,
            in1 => \N__45156\,
            in2 => \_gnd_net_\,
            in3 => \N__36829\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48789\,
            ce => \N__45212\,
            sr => \N__48126\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37005\,
            in2 => \_gnd_net_\,
            in3 => \N__37108\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48781\,
            ce => \N__45211\,
            sr => \N__48130\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__37129\,
            in1 => \_gnd_net_\,
            in2 => \N__37012\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48781\,
            ce => \N__45211\,
            sr => \N__48130\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37009\,
            in2 => \_gnd_net_\,
            in3 => \N__37180\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48781\,
            ce => \N__45211\,
            sr => \N__48130\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37152\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48781\,
            ce => \N__45211\,
            sr => \N__48130\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__45155\,
            in1 => \_gnd_net_\,
            in2 => \N__38917\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48781\,
            ce => \N__45211\,
            sr => \N__48130\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39364\,
            lcout => \current_shift_inst.un4_control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39355\,
            lcout => \current_shift_inst.un4_control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39346\,
            lcout => \current_shift_inst.un4_control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39123\,
            in2 => \_gnd_net_\,
            in3 => \N__46386\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37179\,
            in1 => \N__37128\,
            in2 => \N__37153\,
            in3 => \N__37107\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39337\,
            lcout => \current_shift_inst.un4_control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39328\,
            lcout => \current_shift_inst.un4_control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39319\,
            lcout => \current_shift_inst.un4_control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39310\,
            lcout => \current_shift_inst.un4_control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39301\,
            lcout => \current_shift_inst.un4_control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39493\,
            lcout => \current_shift_inst.un4_control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39292\,
            lcout => \current_shift_inst.un4_control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39382\,
            lcout => \current_shift_inst.un4_control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39400\,
            lcout => \current_shift_inst.un4_control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39418\,
            lcout => \current_shift_inst.un4_control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39409\,
            lcout => \current_shift_inst.un4_control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39391\,
            lcout => \current_shift_inst.un4_control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39484\,
            lcout => \current_shift_inst.un4_control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39454\,
            lcout => \current_shift_inst.un4_control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39373\,
            lcout => \current_shift_inst.un4_control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39889\,
            lcout => \current_shift_inst.un4_control_input_axb_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39463\,
            lcout => \current_shift_inst.un4_control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39898\,
            lcout => \current_shift_inst.un4_control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39445\,
            lcout => \current_shift_inst.un4_control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39472\,
            lcout => \current_shift_inst.un4_control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36989\,
            in2 => \_gnd_net_\,
            in3 => \N__37106\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48750\,
            ce => \N__46643\,
            sr => \N__48154\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37127\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48750\,
            ce => \N__46643\,
            sr => \N__48154\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36991\,
            in2 => \_gnd_net_\,
            in3 => \N__37172\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48750\,
            ce => \N__46643\,
            sr => \N__48154\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37148\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48750\,
            ce => \N__46643\,
            sr => \N__48154\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39502\,
            lcout => \current_shift_inst.un4_control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39433\,
            lcout => \current_shift_inst.un4_control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__49102\,
            in1 => \N__44081\,
            in2 => \_gnd_net_\,
            in3 => \N__46696\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__44082\,
            in1 => \N__49103\,
            in2 => \_gnd_net_\,
            in3 => \N__47482\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__46417\,
            in1 => \N__46502\,
            in2 => \N__45973\,
            in3 => \N__46165\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__44080\,
            in1 => \N__49101\,
            in2 => \_gnd_net_\,
            in3 => \N__46744\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__49100\,
            in1 => \N__44079\,
            in2 => \_gnd_net_\,
            in3 => \N__46789\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010111001111"
        )
    port map (
            in0 => \N__46503\,
            in1 => \N__47020\,
            in2 => \N__46168\,
            in3 => \N__46418\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__44083\,
            in1 => \N__49104\,
            in2 => \N__46864\,
            in3 => \N__46416\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48744\,
            ce => \N__46343\,
            sr => \N__48161\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_2_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40084\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48737\,
            ce => \N__41821\,
            sr => \N__48171\
        );

    \current_shift_inst.un38_control_input_0_cry_3_c_inv_RNO_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100101"
        )
    port map (
            in0 => \N__40101\,
            in1 => \N__37286\,
            in2 => \N__37443\,
            in3 => \N__37321\,
            lcout => \current_shift_inst.N_1742_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_1_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40129\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48737\,
            ce => \N__41821\,
            sr => \N__48171\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_RNI5LGN1_3_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__37322\,
            in1 => \N__40102\,
            in2 => \N__37293\,
            in3 => \N__37431\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5LGN1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_1_c_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37317\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.z_5_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_2_s_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37285\,
            in2 => \N__43357\,
            in3 => \N__37258\,
            lcout => \current_shift_inst.z_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_1\,
            carryout => \current_shift_inst.z_5_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_3_s_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40095\,
            in2 => \N__43361\,
            in3 => \N__37246\,
            lcout => \current_shift_inst.z_5_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_2\,
            carryout => \current_shift_inst.z_5_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_4_s_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40037\,
            in2 => \N__43358\,
            in3 => \N__37231\,
            lcout => \current_shift_inst.z_5_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_3\,
            carryout => \current_shift_inst.z_5_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_5_s_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39971\,
            in2 => \N__43362\,
            in3 => \N__37219\,
            lcout => \current_shift_inst.z_5_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_4\,
            carryout => \current_shift_inst.z_5_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_6_s_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39917\,
            in2 => \N__43359\,
            in3 => \N__37204\,
            lcout => \current_shift_inst.z_5_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_5\,
            carryout => \current_shift_inst.z_5_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_7_s_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40679\,
            in2 => \N__43363\,
            in3 => \N__37567\,
            lcout => \current_shift_inst.z_5_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_6\,
            carryout => \current_shift_inst.z_5_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_8_s_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40606\,
            in2 => \N__43360\,
            in3 => \N__37552\,
            lcout => \current_shift_inst.z_5_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_7\,
            carryout => \current_shift_inst.z_5_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_9_s_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40541\,
            in2 => \N__43467\,
            in3 => \N__37537\,
            lcout => \current_shift_inst.z_5_9\,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \current_shift_inst.z_5_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_10_s_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40472\,
            in2 => \N__43450\,
            in3 => \N__37525\,
            lcout => \current_shift_inst.z_5_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_9\,
            carryout => \current_shift_inst.z_5_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_11_s_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40393\,
            in2 => \N__43464\,
            in3 => \N__37513\,
            lcout => \current_shift_inst.z_5_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_10\,
            carryout => \current_shift_inst.z_5_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_12_s_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40319\,
            in2 => \N__43451\,
            in3 => \N__37498\,
            lcout => \current_shift_inst.z_5_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_11\,
            carryout => \current_shift_inst.z_5_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_13_s_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40243\,
            in2 => \N__43465\,
            in3 => \N__37486\,
            lcout => \current_shift_inst.z_5_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_12\,
            carryout => \current_shift_inst.z_5_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_14_s_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40163\,
            in2 => \N__43452\,
            in3 => \N__37468\,
            lcout => \current_shift_inst.z_5_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_13\,
            carryout => \current_shift_inst.z_5_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_15_s_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41159\,
            in2 => \N__43466\,
            in3 => \N__37690\,
            lcout => \current_shift_inst.z_5_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_14\,
            carryout => \current_shift_inst.z_5_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_16_s_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41090\,
            in2 => \N__43453\,
            in3 => \N__37672\,
            lcout => \current_shift_inst.z_5_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_15\,
            carryout => \current_shift_inst.z_5_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_17_s_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41021\,
            in2 => \N__43454\,
            in3 => \N__37657\,
            lcout => \current_shift_inst.z_5_17\,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \current_shift_inst.z_5_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_18_s_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40958\,
            in2 => \N__43468\,
            in3 => \N__37639\,
            lcout => \current_shift_inst.z_5_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_17\,
            carryout => \current_shift_inst.z_5_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_19_s_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40887\,
            in2 => \N__43455\,
            in3 => \N__37627\,
            lcout => \current_shift_inst.z_5_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_18\,
            carryout => \current_shift_inst.z_5_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_20_s_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40814\,
            in2 => \N__43469\,
            in3 => \N__37612\,
            lcout => \current_shift_inst.z_5_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_19\,
            carryout => \current_shift_inst.z_5_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_21_s_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40748\,
            in2 => \N__43456\,
            in3 => \N__37600\,
            lcout => \current_shift_inst.z_5_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_20\,
            carryout => \current_shift_inst.z_5_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_22_s_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41705\,
            in2 => \N__43470\,
            in3 => \N__37585\,
            lcout => \current_shift_inst.z_5_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_21\,
            carryout => \current_shift_inst.z_5_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_23_s_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41638\,
            in2 => \N__43457\,
            in3 => \N__37840\,
            lcout => \current_shift_inst.z_5_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_22\,
            carryout => \current_shift_inst.z_5_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_24_s_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41570\,
            in2 => \N__43471\,
            in3 => \N__37822\,
            lcout => \current_shift_inst.z_5_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_23\,
            carryout => \current_shift_inst.z_5_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_25_s_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41510\,
            in2 => \N__43458\,
            in3 => \N__37807\,
            lcout => \current_shift_inst.z_5_25\,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \current_shift_inst.z_5_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_26_s_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41450\,
            in2 => \N__43461\,
            in3 => \N__37789\,
            lcout => \current_shift_inst.z_5_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_25\,
            carryout => \current_shift_inst.z_5_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_27_s_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41384\,
            in2 => \N__43459\,
            in3 => \N__37771\,
            lcout => \current_shift_inst.z_5_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_26\,
            carryout => \current_shift_inst.z_5_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_28_s_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41311\,
            in2 => \N__43462\,
            in3 => \N__37756\,
            lcout => \current_shift_inst.z_5_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_27\,
            carryout => \current_shift_inst.z_5_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_29_s_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41231\,
            in2 => \N__43460\,
            in3 => \N__37738\,
            lcout => \current_shift_inst.z_5_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_28\,
            carryout => \current_shift_inst.z_5_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_z_5_cry_30_s_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41873\,
            in2 => \N__43463\,
            in3 => \N__37723\,
            lcout => \current_shift_inst.z_5_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.z_5_cry_29\,
            carryout => \current_shift_inst.z_5_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.z_5_cry_30_THRU_LUT4_0_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37720\,
            lcout => \current_shift_inst.z_5_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC1_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48862\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37957\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37948\,
            in2 => \N__37942\,
            in3 => \N__44393\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37924\,
            in2 => \N__37933\,
            in3 => \N__44376\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44340\,
            in1 => \N__37909\,
            in2 => \N__37918\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37891\,
            in2 => \N__37903\,
            in3 => \N__44319\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37876\,
            in2 => \N__37885\,
            in3 => \N__44292\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37861\,
            in2 => \N__37870\,
            in3 => \N__44268\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44244\,
            in1 => \N__38098\,
            in2 => \N__38110\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44748\,
            in1 => \N__38083\,
            in2 => \N__38092\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38068\,
            in2 => \N__38077\,
            in3 => \N__44721\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44694\,
            in1 => \N__38053\,
            in2 => \N__38062\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38038\,
            in2 => \N__38047\,
            in3 => \N__44673\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38020\,
            in2 => \N__38032\,
            in3 => \N__44652\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38005\,
            in2 => \N__38014\,
            in3 => \N__44631\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37981\,
            in2 => \N__37999\,
            in3 => \N__44610\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38194\,
            in2 => \N__38206\,
            in3 => \N__44589\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38176\,
            in2 => \N__38188\,
            in3 => \N__44943\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38158\,
            in2 => \N__38170\,
            in3 => \N__44922\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__44889\,
            in1 => \N__38140\,
            in2 => \N__38152\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38119\,
            in2 => \N__38134\,
            in3 => \N__44865\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38113\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42630\,
            in2 => \_gnd_net_\,
            in3 => \N__42590\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__42591\,
            in1 => \_gnd_net_\,
            in2 => \N__42634\,
            in3 => \N__44397\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38386\,
            in2 => \N__39244\,
            in3 => \N__38402\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38379\,
            in1 => \N__38368\,
            in2 => \N__39058\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38358\,
            in1 => \N__38347\,
            in2 => \N__39232\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38317\,
            in2 => \N__38341\,
            in3 => \N__38328\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38299\,
            in2 => \N__38758\,
            in3 => \N__38310\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38269\,
            in2 => \N__38293\,
            in3 => \N__38280\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38239\,
            in2 => \N__38263\,
            in3 => \N__38250\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38626\,
            in2 => \N__38233\,
            in3 => \N__38217\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38599\,
            in2 => \N__38620\,
            in3 => \N__38610\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38560\,
            in2 => \N__38593\,
            in3 => \N__38577\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38542\,
            in2 => \N__38554\,
            in3 => \N__45774\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38512\,
            in2 => \N__38536\,
            in3 => \N__38523\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38502\,
            in1 => \N__38476\,
            in2 => \N__38491\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38446\,
            in2 => \N__38470\,
            in3 => \N__38457\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38413\,
            in2 => \N__38440\,
            in3 => \N__38424\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45235\,
            in2 => \N__38722\,
            in3 => \N__38733\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38701\,
            in2 => \N__38653\,
            in3 => \N__38712\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38680\,
            in2 => \N__38644\,
            in3 => \N__38691\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38662\,
            in2 => \N__38635\,
            in3 => \N__38673\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38656\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39787\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48798\,
            ce => \N__45223\,
            sr => \N__48121\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39831\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48798\,
            ce => \N__45223\,
            sr => \N__48121\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39741\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48798\,
            ce => \N__45223\,
            sr => \N__48121\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__39279\,
            in1 => \N__39146\,
            in2 => \N__39268\,
            in3 => \N__39089\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => \N__45219\,
            sr => \N__48127\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__39091\,
            in1 => \_gnd_net_\,
            in2 => \N__39150\,
            in3 => \N__39129\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => \N__45219\,
            sr => \N__48127\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__38824\,
            in1 => \N__39215\,
            in2 => \N__38926\,
            in3 => \N__39181\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__39130\,
            in1 => \N__46390\,
            in2 => \N__39094\,
            in3 => \N__39090\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => \N__45219\,
            sr => \N__48127\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_6_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__39046\,
            in1 => \N__39002\,
            in2 => \_gnd_net_\,
            in3 => \N__38954\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38913\,
            in2 => \N__38836\,
            in3 => \N__38823\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__38800\,
            in1 => \N__45141\,
            in2 => \N__38761\,
            in3 => \N__44975\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48790\,
            ce => \N__45219\,
            sr => \N__48127\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42498\,
            in2 => \N__42567\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42474\,
            in2 => \N__42531\,
            in3 => \N__39358\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42499\,
            in2 => \N__42450\,
            in3 => \N__39349\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42475\,
            in2 => \N__42420\,
            in3 => \N__39340\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42390\,
            in2 => \N__42451\,
            in3 => \N__39331\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42366\,
            in2 => \N__42421\,
            in3 => \N__39322\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42391\,
            in2 => \N__42859\,
            in3 => \N__39313\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42367\,
            in2 => \N__42828\,
            in3 => \N__39304\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__48782\,
            ce => \N__39880\,
            sr => \N__48131\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42858\,
            in2 => \N__42796\,
            in3 => \N__39295\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42765\,
            in2 => \N__42829\,
            in3 => \N__39436\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42795\,
            in2 => \N__42741\,
            in3 => \N__39424\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42766\,
            in2 => \N__42711\,
            in3 => \N__39421\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42681\,
            in2 => \N__42742\,
            in3 => \N__39412\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42657\,
            in2 => \N__42712\,
            in3 => \N__39403\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42682\,
            in2 => \N__43114\,
            in3 => \N__39394\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42658\,
            in2 => \N__43084\,
            in3 => \N__39385\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__48773\,
            ce => \N__39879\,
            sr => \N__48136\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43113\,
            in2 => \N__43053\,
            in3 => \N__39376\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_16_17_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43083\,
            in2 => \N__43024\,
            in3 => \N__39367\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42993\,
            in2 => \N__43054\,
            in3 => \N__39496\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43023\,
            in2 => \N__42969\,
            in3 => \N__39487\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42994\,
            in2 => \N__42940\,
            in3 => \N__39478\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42909\,
            in2 => \N__42970\,
            in3 => \N__39475\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42939\,
            in2 => \N__42886\,
            in3 => \N__39466\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42910\,
            in2 => \N__43837\,
            in3 => \N__39457\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__48763\,
            ce => \N__39877\,
            sr => \N__48142\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42885\,
            in2 => \N__43806\,
            in3 => \N__39448\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__48756\,
            ce => \N__39876\,
            sr => \N__48148\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43836\,
            in2 => \N__43777\,
            in3 => \N__39439\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__48756\,
            ce => \N__39876\,
            sr => \N__48148\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43747\,
            in2 => \N__43807\,
            in3 => \N__39892\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__48756\,
            ce => \N__39876\,
            sr => \N__48148\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43776\,
            in2 => \N__43597\,
            in3 => \N__39883\,
            lcout => \current_shift_inst.timer_s1.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__48756\,
            ce => \N__39876\,
            sr => \N__48148\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39856\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__39824\,
            in1 => \N__39782\,
            in2 => \N__39745\,
            in3 => \N__45263\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5PP_2_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__46474\,
            in1 => \N__47428\,
            in2 => \N__46086\,
            in3 => \N__46030\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__46916\,
            in1 => \N__46970\,
            in2 => \_gnd_net_\,
            in3 => \N__47019\,
            lcout => \delay_measurement_inst.N_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.T01_sbtinv_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__39690\,
            in1 => \N__39642\,
            in2 => \N__39604\,
            in3 => \N__39553\,
            lcout => \phase_controller_inst1.N_221_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9DQM6_10_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44097\,
            in2 => \_gnd_net_\,
            in3 => \N__46219\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_424_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__40147\,
            in1 => \N__46501\,
            in2 => \N__39505\,
            in3 => \N__40138\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__47354\,
            in1 => \N__44098\,
            in2 => \_gnd_net_\,
            in3 => \N__46220\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI86841_4_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47418\,
            in1 => \N__46029\,
            in2 => \N__47363\,
            in3 => \N__45968\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICTS5M_31_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48275\,
            in2 => \_gnd_net_\,
            in3 => \N__43851\,
            lcout => \delay_measurement_inst.N_280_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47172\,
            in1 => \N__47232\,
            in2 => \N__47117\,
            in3 => \N__47289\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__46079\,
            in1 => \N__46463\,
            in2 => \N__40141\,
            in3 => \N__46852\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_3_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40125\,
            in2 => \N__40018\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_3\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_4_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40082\,
            in2 => \N__39955\,
            in3 => \N__40021\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_5_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40017\,
            in2 => \N__40728\,
            in3 => \N__39958\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_6_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39954\,
            in2 => \N__40659\,
            in3 => \N__39901\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_7_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40581\,
            in2 => \N__40729\,
            in3 => \N__40663\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_8_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40521\,
            in2 => \N__40660\,
            in3 => \N__40585\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_9_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40582\,
            in2 => \N__40453\,
            in3 => \N__40525\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_10_LC_16_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40522\,
            in2 => \N__40369\,
            in3 => \N__40456\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_9\,
            clk => \N__48732\,
            ce => \N__41820\,
            sr => \N__48184\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_11_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40446\,
            in2 => \N__40299\,
            in3 => \N__40372\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_11\,
            ltout => OPEN,
            carryin => \bfn_16_23_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_12_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40368\,
            in2 => \N__40219\,
            in3 => \N__40303\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_13_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41208\,
            in2 => \N__40300\,
            in3 => \N__40222\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_14_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40218\,
            in2 => \N__41139\,
            in3 => \N__41212\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_15_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41209\,
            in2 => \N__41070\,
            in3 => \N__41143\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_16_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41001\,
            in2 => \N__41140\,
            in3 => \N__41074\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_17_LC_16_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40939\,
            in2 => \N__41071\,
            in3 => \N__41005\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_18_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41002\,
            in2 => \N__40873\,
            in3 => \N__40942\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_17\,
            clk => \N__48725\,
            ce => \N__41819\,
            sr => \N__48192\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_19_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40938\,
            in2 => \N__40795\,
            in3 => \N__40876\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_19\,
            ltout => OPEN,
            carryin => \bfn_16_24_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_20_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40866\,
            in2 => \N__41752\,
            in3 => \N__40798\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_21_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40794\,
            in2 => \N__41685\,
            in3 => \N__40732\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_22_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41751\,
            in2 => \N__41613\,
            in3 => \N__41689\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_23_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41547\,
            in2 => \N__41686\,
            in3 => \N__41617\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_24_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41490\,
            in2 => \N__41614\,
            in3 => \N__41554\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_25_LC_16_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41431\,
            in2 => \N__41551\,
            in3 => \N__41494\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_26_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41491\,
            in2 => \N__41365\,
            in3 => \N__41434\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_25\,
            clk => \N__48718\,
            ce => \N__41818\,
            sr => \N__48199\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_27_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41430\,
            in2 => \N__41271\,
            in3 => \N__41368\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_27\,
            ltout => OPEN,
            carryin => \bfn_16_25_0_\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            clk => \N__48712\,
            ce => \N__41817\,
            sr => \N__48207\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_28_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41364\,
            in2 => \N__41932\,
            in3 => \N__41290\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            clk => \N__48712\,
            ce => \N__41817\,
            sr => \N__48207\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_29_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41287\,
            in2 => \N__41272\,
            in3 => \N__41215\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            clk => \N__48712\,
            ce => \N__41817\,
            sr => \N__48207\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_30_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41931\,
            in2 => \N__41908\,
            in3 => \N__41857\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_phase.un13_elapsed_time_ns_cry_29\,
            clk => \N__48712\,
            ce => \N__41817\,
            sr => \N__48207\
        );

    \current_shift_inst.timer_phase.elapsed_time_ns_1_31_LC_16_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41854\,
            lcout => \current_shift_inst.elapsed_time_ns_phase_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48712\,
            ce => \N__41817\,
            sr => \N__48207\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_16_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47548\,
            in1 => \N__47581\,
            in2 => \N__47518\,
            in3 => \N__47617\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47056\,
            in1 => \N__41797\,
            in2 => \N__41800\,
            in3 => \N__41791\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__47686\,
            in1 => \N__47716\,
            in2 => \N__47656\,
            in3 => \N__47752\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO4MS_29_LC_16_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49144\,
            in2 => \_gnd_net_\,
            in3 => \N__49192\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41782\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41767\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42310\,
            in1 => \N__42174\,
            in2 => \N__44281\,
            in3 => \N__42057\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42054\,
            in1 => \N__42314\,
            in2 => \N__42190\,
            in3 => \N__44737\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42308\,
            in1 => \N__42172\,
            in2 => \N__44905\,
            in3 => \N__42055\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42051\,
            in1 => \N__42311\,
            in2 => \N__42187\,
            in3 => \N__44365\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42053\,
            in1 => \N__42313\,
            in2 => \N__42189\,
            in3 => \N__44257\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__42309\,
            in1 => \N__42173\,
            in2 => \N__44308\,
            in3 => \N__42056\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42052\,
            in1 => \N__42312\,
            in2 => \N__42188\,
            in3 => \N__44329\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48847\,
            ce => 'H',
            sr => \N__48088\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__42315\,
            in1 => \N__42047\,
            in2 => \N__42175\,
            in3 => \N__44683\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42045\,
            in1 => \N__42136\,
            in2 => \N__42333\,
            in3 => \N__44878\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__42317\,
            in1 => \N__42049\,
            in2 => \N__42177\,
            in3 => \N__44641\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42043\,
            in1 => \N__42134\,
            in2 => \N__42331\,
            in3 => \N__44620\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__42318\,
            in1 => \N__42050\,
            in2 => \N__42178\,
            in3 => \N__44578\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42044\,
            in1 => \N__42135\,
            in2 => \N__42332\,
            in3 => \N__44599\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__42316\,
            in1 => \N__42048\,
            in2 => \N__42176\,
            in3 => \N__44662\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__42046\,
            in1 => \N__42137\,
            in2 => \N__42334\,
            in3 => \N__42343\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48841\,
            ce => 'H',
            sr => \N__48090\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44798\,
            in2 => \_gnd_net_\,
            in3 => \N__44821\,
            lcout => OPEN,
            ltout => \phase_controller_slave.N_214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__42132\,
            in1 => \N__44833\,
            in2 => \N__42337\,
            in3 => \N__45937\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48836\,
            ce => 'H',
            sr => \N__48093\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__42305\,
            in1 => \N__42133\,
            in2 => \N__42061\,
            in3 => \N__44932\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48836\,
            ce => 'H',
            sr => \N__48093\
        );

    \phase_controller_slave.state_2_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__44822\,
            in1 => \N__45822\,
            in2 => \N__44805\,
            in3 => \N__45760\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48836\,
            ce => 'H',
            sr => \N__48093\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__44823\,
            in1 => \N__42629\,
            in2 => \N__41944\,
            in3 => \N__42589\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48836\,
            ce => 'H',
            sr => \N__48093\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42628\,
            in2 => \_gnd_net_\,
            in3 => \N__42588\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43703\,
            in1 => \N__42554\,
            in2 => \_gnd_net_\,
            in3 => \N__42538\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43711\,
            in1 => \N__42518\,
            in2 => \_gnd_net_\,
            in3 => \N__42502\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43704\,
            in1 => \N__42497\,
            in2 => \_gnd_net_\,
            in3 => \N__42478\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_3_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43712\,
            in1 => \N__42468\,
            in2 => \_gnd_net_\,
            in3 => \N__42454\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_4_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43705\,
            in1 => \N__42438\,
            in2 => \_gnd_net_\,
            in3 => \N__42424\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_5_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43713\,
            in1 => \N__42408\,
            in2 => \_gnd_net_\,
            in3 => \N__42394\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_6_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43706\,
            in1 => \N__42384\,
            in2 => \_gnd_net_\,
            in3 => \N__42370\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_7_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43714\,
            in1 => \N__42360\,
            in2 => \_gnd_net_\,
            in3 => \N__42346\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__48827\,
            ce => \N__43576\,
            sr => \N__48099\
        );

    \current_shift_inst.timer_s1.counter_8_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43718\,
            in1 => \N__42848\,
            in2 => \_gnd_net_\,
            in3 => \N__42832\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_9_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43726\,
            in1 => \N__42815\,
            in2 => \_gnd_net_\,
            in3 => \N__42799\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_10_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43715\,
            in1 => \N__42791\,
            in2 => \_gnd_net_\,
            in3 => \N__42769\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_11_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43723\,
            in1 => \N__42764\,
            in2 => \_gnd_net_\,
            in3 => \N__42745\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_12_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43716\,
            in1 => \N__42729\,
            in2 => \_gnd_net_\,
            in3 => \N__42715\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_13_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43724\,
            in1 => \N__42699\,
            in2 => \_gnd_net_\,
            in3 => \N__42685\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_14_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43717\,
            in1 => \N__42675\,
            in2 => \_gnd_net_\,
            in3 => \N__42661\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_15_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43725\,
            in1 => \N__42651\,
            in2 => \_gnd_net_\,
            in3 => \N__42637\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__48817\,
            ce => \N__43571\,
            sr => \N__48107\
        );

    \current_shift_inst.timer_s1.counter_16_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43707\,
            in1 => \N__43103\,
            in2 => \_gnd_net_\,
            in3 => \N__43087\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_17_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43719\,
            in1 => \N__43073\,
            in2 => \_gnd_net_\,
            in3 => \N__43057\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_18_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43708\,
            in1 => \N__43046\,
            in2 => \_gnd_net_\,
            in3 => \N__43027\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_19_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43720\,
            in1 => \N__43019\,
            in2 => \_gnd_net_\,
            in3 => \N__42997\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_20_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43709\,
            in1 => \N__42987\,
            in2 => \_gnd_net_\,
            in3 => \N__42973\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_21_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43721\,
            in1 => \N__42957\,
            in2 => \_gnd_net_\,
            in3 => \N__42943\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_22_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43710\,
            in1 => \N__42929\,
            in2 => \_gnd_net_\,
            in3 => \N__42913\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_23_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43722\,
            in1 => \N__42903\,
            in2 => \_gnd_net_\,
            in3 => \N__42889\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__48810\,
            ce => \N__43561\,
            sr => \N__48113\
        );

    \current_shift_inst.timer_s1.counter_24_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43643\,
            in1 => \N__42875\,
            in2 => \_gnd_net_\,
            in3 => \N__43840\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_14_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__48799\,
            ce => \N__43572\,
            sr => \N__48122\
        );

    \current_shift_inst.timer_s1.counter_25_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43647\,
            in1 => \N__43826\,
            in2 => \_gnd_net_\,
            in3 => \N__43810\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__48799\,
            ce => \N__43572\,
            sr => \N__48122\
        );

    \current_shift_inst.timer_s1.counter_26_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43644\,
            in1 => \N__43799\,
            in2 => \_gnd_net_\,
            in3 => \N__43780\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__48799\,
            ce => \N__43572\,
            sr => \N__48122\
        );

    \current_shift_inst.timer_s1.counter_27_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43648\,
            in1 => \N__43772\,
            in2 => \_gnd_net_\,
            in3 => \N__43750\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__48799\,
            ce => \N__43572\,
            sr => \N__48122\
        );

    \current_shift_inst.timer_s1.counter_28_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__43645\,
            in1 => \N__43743\,
            in2 => \_gnd_net_\,
            in3 => \N__43729\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__48799\,
            ce => \N__43572\,
            sr => \N__48122\
        );

    \current_shift_inst.timer_s1.counter_29_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__43590\,
            in1 => \N__43646\,
            in2 => \_gnd_net_\,
            in3 => \N__43600\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48799\,
            ce => \N__43572\,
            sr => \N__48122\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43531\,
            lcout => \current_shift_inst.un4_control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43516\,
            lcout => \current_shift_inst.un4_control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_tr_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43985\,
            in1 => \N__44014\,
            in2 => \_gnd_net_\,
            in3 => \N__43943\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48143\
        );

    \delay_measurement_inst.prev_tr_sig_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43986\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48143\
        );

    \delay_measurement_inst.stop_timer_tr_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43908\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48143\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__44131\,
            in1 => \N__44116\,
            in2 => \_gnd_net_\,
            in3 => \N__44058\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48764\,
            ce => 'H',
            sr => \N__48143\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9IAF_1_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__47018\,
            in1 => \N__45969\,
            in2 => \N__46860\,
            in3 => \N__48895\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI200N_7_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__46917\,
            in1 => \_gnd_net_\,
            in2 => \N__43924\,
            in3 => \N__46971\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_2_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__43921\,
            in1 => \N__46268\,
            in2 => \N__43915\,
            in3 => \N__46415\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.N_390_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5KUTL_31_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__49095\,
            in1 => \N__43912\,
            in2 => \N__43888\,
            in3 => \N__43885\,
            lcout => \delay_measurement_inst.N_280_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44114\,
            in2 => \_gnd_net_\,
            in3 => \N__44056\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_338_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__44057\,
            in1 => \N__44127\,
            in2 => \_gnd_net_\,
            in3 => \N__44115\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_339_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46692\,
            in1 => \N__46740\,
            in2 => \N__47481\,
            in3 => \N__46788\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110001"
        )
    port map (
            in0 => \N__47425\,
            in1 => \N__47361\,
            in2 => \N__44086\,
            in3 => \N__46856\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001101"
        )
    port map (
            in0 => \N__47426\,
            in1 => \N__46270\,
            in2 => \N__47364\,
            in3 => \N__46241\,
            lcout => \delay_measurement_inst.N_409_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44059\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46051\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48745\,
            ce => \N__48338\,
            sr => \N__48162\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45270\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48738\,
            ce => \N__46648\,
            sr => \N__48172\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44545\,
            in1 => \N__48911\,
            in2 => \_gnd_net_\,
            in3 => \N__44020\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44540\,
            in1 => \N__46046\,
            in2 => \_gnd_net_\,
            in3 => \N__44017\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44546\,
            in1 => \N__45992\,
            in2 => \_gnd_net_\,
            in3 => \N__44158\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44541\,
            in1 => \N__47039\,
            in2 => \_gnd_net_\,
            in3 => \N__44155\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44547\,
            in1 => \N__46993\,
            in2 => \_gnd_net_\,
            in3 => \N__44152\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44542\,
            in1 => \N__46939\,
            in2 => \_gnd_net_\,
            in3 => \N__44149\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44544\,
            in1 => \N__46883\,
            in2 => \_gnd_net_\,
            in3 => \N__44146\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44543\,
            in1 => \N__46808\,
            in2 => \_gnd_net_\,
            in3 => \N__44143\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__48733\,
            ce => \N__44440\,
            sr => \N__48185\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44551\,
            in1 => \N__46761\,
            in2 => \_gnd_net_\,
            in3 => \N__44140\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44569\,
            in1 => \N__46713\,
            in2 => \_gnd_net_\,
            in3 => \N__44137\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44548\,
            in1 => \N__47501\,
            in2 => \_gnd_net_\,
            in3 => \N__44134\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44566\,
            in1 => \N__47447\,
            in2 => \_gnd_net_\,
            in3 => \N__44185\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44549\,
            in1 => \N__47380\,
            in2 => \_gnd_net_\,
            in3 => \N__44182\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44567\,
            in1 => \N__47308\,
            in2 => \_gnd_net_\,
            in3 => \N__44179\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44550\,
            in1 => \N__47252\,
            in2 => \_gnd_net_\,
            in3 => \N__44176\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44568\,
            in1 => \N__47198\,
            in2 => \_gnd_net_\,
            in3 => \N__44173\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__48726\,
            ce => \N__44442\,
            sr => \N__48193\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44552\,
            in1 => \N__47139\,
            in2 => \_gnd_net_\,
            in3 => \N__44170\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_25_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44556\,
            in1 => \N__47073\,
            in2 => \_gnd_net_\,
            in3 => \N__44167\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44553\,
            in1 => \N__47771\,
            in2 => \_gnd_net_\,
            in3 => \N__44164\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44557\,
            in1 => \N__47735\,
            in2 => \_gnd_net_\,
            in3 => \N__44161\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44554\,
            in1 => \N__47701\,
            in2 => \_gnd_net_\,
            in3 => \N__44212\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44558\,
            in1 => \N__47671\,
            in2 => \_gnd_net_\,
            in3 => \N__44209\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44555\,
            in1 => \N__47636\,
            in2 => \_gnd_net_\,
            in3 => \N__44206\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44559\,
            in1 => \N__47600\,
            in2 => \_gnd_net_\,
            in3 => \N__44203\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__48719\,
            ce => \N__44441\,
            sr => \N__48200\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44560\,
            in1 => \N__47565\,
            in2 => \_gnd_net_\,
            in3 => \N__44200\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__48713\,
            ce => \N__44443\,
            sr => \N__48208\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44564\,
            in1 => \N__47535\,
            in2 => \_gnd_net_\,
            in3 => \N__44197\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__48713\,
            ce => \N__44443\,
            sr => \N__48208\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44561\,
            in1 => \N__49211\,
            in2 => \_gnd_net_\,
            in3 => \N__44194\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__48713\,
            ce => \N__44443\,
            sr => \N__48208\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44565\,
            in1 => \N__49163\,
            in2 => \_gnd_net_\,
            in3 => \N__44191\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__48713\,
            ce => \N__44443\,
            sr => \N__48208\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44562\,
            in1 => \N__49225\,
            in2 => \_gnd_net_\,
            in3 => \N__44188\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__48713\,
            ce => \N__44443\,
            sr => \N__48208\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__49177\,
            in1 => \N__44563\,
            in2 => \_gnd_net_\,
            in3 => \N__44446\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48713\,
            ce => \N__44443\,
            sr => \N__48208\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44407\,
            in2 => \N__44398\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_8_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44377\,
            in2 => \_gnd_net_\,
            in3 => \N__44359\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44356\,
            in2 => \N__44344\,
            in3 => \N__44323\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44320\,
            in2 => \_gnd_net_\,
            in3 => \N__44296\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44293\,
            in2 => \_gnd_net_\,
            in3 => \N__44272\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44269\,
            in2 => \_gnd_net_\,
            in3 => \N__44251\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44248\,
            in2 => \_gnd_net_\,
            in3 => \N__44215\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44749\,
            in2 => \_gnd_net_\,
            in3 => \N__44731\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44728\,
            in2 => \_gnd_net_\,
            in3 => \N__44698\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_18_9_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44695\,
            in2 => \_gnd_net_\,
            in3 => \N__44677\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44674\,
            in2 => \_gnd_net_\,
            in3 => \N__44656\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44653\,
            in2 => \_gnd_net_\,
            in3 => \N__44635\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44632\,
            in2 => \_gnd_net_\,
            in3 => \N__44614\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44611\,
            in2 => \_gnd_net_\,
            in3 => \N__44593\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44590\,
            in2 => \_gnd_net_\,
            in3 => \N__44572\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44944\,
            in2 => \_gnd_net_\,
            in3 => \N__44926\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44923\,
            in2 => \_gnd_net_\,
            in3 => \N__44893\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_18_10_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44890\,
            in2 => \_gnd_net_\,
            in3 => \N__44872\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44869\,
            in2 => \_gnd_net_\,
            in3 => \N__44848\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45759\,
            in2 => \_gnd_net_\,
            in3 => \N__45818\,
            lcout => \phase_controller_slave.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_1_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__44824\,
            in1 => \N__49035\,
            in2 => \N__44806\,
            in3 => \N__49013\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48837\,
            ce => 'H',
            sr => \N__48094\
        );

    \phase_controller_slave.S2_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__45757\,
            in1 => \N__49034\,
            in2 => \N__44766\,
            in3 => \N__45727\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48837\,
            ce => 'H',
            sr => \N__48094\
        );

    \phase_controller_slave.state_0_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__49014\,
            in1 => \N__48971\,
            in2 => \N__49039\,
            in3 => \N__48948\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48837\,
            ce => 'H',
            sr => \N__48094\
        );

    \phase_controller_slave.start_timer_tr_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__48985\,
            in1 => \N__45930\,
            in2 => \N__45603\,
            in3 => \N__48934\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48828\,
            ce => 'H',
            sr => \N__48100\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__45555\,
            in1 => \N__45460\,
            in2 => \_gnd_net_\,
            in3 => \N__45392\,
            lcout => OPEN,
            ltout => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__48972\,
            in1 => \N__45904\,
            in2 => \N__45877\,
            in3 => \N__45874\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48828\,
            ce => 'H',
            sr => \N__48100\
        );

    \phase_controller_slave.state_3_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__48933\,
            in1 => \N__45758\,
            in2 => \N__45823\,
            in3 => \N__45796\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48828\,
            ce => 'H',
            sr => \N__48100\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__45393\,
            in1 => \N__45556\,
            in2 => \N__45498\,
            in3 => \N__45787\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48828\,
            ce => 'H',
            sr => \N__48100\
        );

    \phase_controller_slave.S1_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__45666\,
            in1 => \N__45756\,
            in2 => \_gnd_net_\,
            in3 => \N__45726\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48818\,
            ce => 'H',
            sr => \N__48108\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__45560\,
            in1 => \N__45459\,
            in2 => \_gnd_net_\,
            in3 => \N__45326\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45274\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48800\,
            ce => \N__45196\,
            sr => \N__48123\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__45137\,
            in1 => \N__45052\,
            in2 => \N__46559\,
            in3 => \N__44993\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48783\,
            ce => \N__46644\,
            sr => \N__48132\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__46028\,
            in1 => \N__46526\,
            in2 => \N__46153\,
            in3 => \N__46439\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48774\,
            ce => \N__46349\,
            sr => \N__48137\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__46516\,
            in1 => \N__46473\,
            in2 => \N__46135\,
            in3 => \N__46438\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48765\,
            ce => \N__46344\,
            sr => \N__48144\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL5GJ7_15_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__47362\,
            in1 => \N__46269\,
            in2 => \N__49114\,
            in3 => \N__46251\,
            lcout => \delay_measurement_inst.N_286_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__47168\,
            in1 => \N__47228\,
            in2 => \N__47118\,
            in3 => \N__47282\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__46252\,
            in1 => \N__49099\,
            in2 => \N__46177\,
            in3 => \N__46174\,
            lcout => \delay_measurement_inst.N_373\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48912\,
            in2 => \N__45993\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_18_23_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46047\,
            in2 => \N__47040\,
            in3 => \N__45997\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46991\,
            in2 => \N__45994\,
            in3 => \N__45940\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46937\,
            in2 => \N__47041\,
            in3 => \N__46996\,
            lcout => \delay_measurement_inst.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46992\,
            in2 => \N__46884\,
            in3 => \N__46942\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46938\,
            in2 => \N__46809\,
            in3 => \N__46888\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46760\,
            in2 => \N__46885\,
            in3 => \N__46813\,
            lcout => \delay_measurement_inst.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46712\,
            in2 => \N__46810\,
            in3 => \N__46765\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__48739\,
            ce => \N__48346\,
            sr => \N__48173\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46762\,
            in2 => \N__47502\,
            in3 => \N__46717\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_18_24_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46714\,
            in2 => \N__47448\,
            in3 => \N__46669\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47378\,
            in2 => \N__47503\,
            in3 => \N__47452\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47306\,
            in2 => \N__47449\,
            in3 => \N__47383\,
            lcout => \delay_measurement_inst.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47379\,
            in2 => \N__47253\,
            in3 => \N__47311\,
            lcout => \delay_measurement_inst.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47307\,
            in2 => \N__47199\,
            in3 => \N__47257\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_18_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47138\,
            in2 => \N__47254\,
            in3 => \N__47203\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47072\,
            in2 => \N__47200\,
            in3 => \N__47143\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__48734\,
            ce => \N__48343\,
            sr => \N__48186\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47140\,
            in2 => \N__47772\,
            in3 => \N__47077\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_18_25_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47074\,
            in2 => \N__47736\,
            in3 => \N__47044\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47699\,
            in2 => \N__47773\,
            in3 => \N__47740\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47669\,
            in2 => \N__47737\,
            in3 => \N__47704\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47700\,
            in2 => \N__47637\,
            in3 => \N__47674\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47670\,
            in2 => \N__47601\,
            in3 => \N__47641\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47564\,
            in2 => \N__47638\,
            in3 => \N__47605\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47534\,
            in2 => \N__47602\,
            in3 => \N__47569\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__48727\,
            ce => \N__48345\,
            sr => \N__48194\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47566\,
            in2 => \N__49212\,
            in3 => \N__47539\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_18_26_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__48720\,
            ce => \N__48344\,
            sr => \N__48201\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47536\,
            in2 => \N__49164\,
            in3 => \N__47506\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__48720\,
            ce => \N__48344\,
            sr => \N__48201\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49224\,
            in2 => \N__49213\,
            in3 => \N__49180\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__48720\,
            ce => \N__48344\,
            sr => \N__48201\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49176\,
            in2 => \N__49165\,
            in3 => \N__49132\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__48720\,
            ce => \N__48344\,
            sr => \N__48201\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49129\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48720\,
            ce => \N__48344\,
            sr => \N__48201\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49033\,
            in2 => \_gnd_net_\,
            in3 => \N__49015\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_RNIVDE2_0_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48973\,
            in2 => \_gnd_net_\,
            in3 => \N__48952\,
            lcout => \phase_controller_slave.N_211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48922\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__48791\,
            ce => \N__48339\,
            sr => \N__48138\
        );
end \INTERFACE\;
