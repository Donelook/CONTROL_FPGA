-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 13 2025 23:22:37

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    rgb_g : out std_logic;
    T01 : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    T23 : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    clock_output : out std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    T45 : out std_logic;
    T12 : out std_logic;
    s4_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48637\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48609\ : std_logic;
signal \N__48608\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48599\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48573\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48555\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48547\ : std_logic;
signal \N__48546\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48538\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48536\ : std_logic;
signal \N__48529\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48500\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48465\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48463\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48449\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48436\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48400\ : std_logic;
signal \N__48397\ : std_logic;
signal \N__48394\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48377\ : std_logic;
signal \N__48376\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48367\ : std_logic;
signal \N__48362\ : std_logic;
signal \N__48359\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48342\ : std_logic;
signal \N__48341\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48339\ : std_logic;
signal \N__48338\ : std_logic;
signal \N__48337\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48334\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48331\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48328\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48309\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48306\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48300\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48298\ : std_logic;
signal \N__48297\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48295\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48289\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48279\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48268\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48260\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48249\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48231\ : std_logic;
signal \N__48230\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48201\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48193\ : std_logic;
signal \N__48192\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48189\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48163\ : std_logic;
signal \N__48152\ : std_logic;
signal \N__48143\ : std_logic;
signal \N__48138\ : std_logic;
signal \N__48135\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48121\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48119\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48115\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48078\ : std_logic;
signal \N__48075\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48073\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48034\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48026\ : std_logic;
signal \N__48019\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48004\ : std_logic;
signal \N__47999\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47971\ : std_logic;
signal \N__47966\ : std_logic;
signal \N__47957\ : std_logic;
signal \N__47954\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47944\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47891\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47841\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47805\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47793\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47777\ : std_logic;
signal \N__47770\ : std_logic;
signal \N__47761\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47735\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47717\ : std_logic;
signal \N__47714\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47671\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47656\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47635\ : std_logic;
signal \N__47632\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47583\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47577\ : std_logic;
signal \N__47576\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47570\ : std_logic;
signal \N__47567\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47555\ : std_logic;
signal \N__47554\ : std_logic;
signal \N__47553\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47551\ : std_logic;
signal \N__47550\ : std_logic;
signal \N__47549\ : std_logic;
signal \N__47548\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47544\ : std_logic;
signal \N__47543\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47541\ : std_logic;
signal \N__47540\ : std_logic;
signal \N__47539\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47537\ : std_logic;
signal \N__47536\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47534\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47531\ : std_logic;
signal \N__47530\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47528\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47525\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47522\ : std_logic;
signal \N__47521\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47519\ : std_logic;
signal \N__47518\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47516\ : std_logic;
signal \N__47515\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47513\ : std_logic;
signal \N__47512\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47506\ : std_logic;
signal \N__47505\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47502\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47500\ : std_logic;
signal \N__47499\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47497\ : std_logic;
signal \N__47496\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47494\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47492\ : std_logic;
signal \N__47491\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47489\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47486\ : std_logic;
signal \N__47485\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47483\ : std_logic;
signal \N__47482\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47480\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47477\ : std_logic;
signal \N__47476\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47474\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47471\ : std_logic;
signal \N__47470\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47467\ : std_logic;
signal \N__47466\ : std_logic;
signal \N__47465\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47462\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47459\ : std_logic;
signal \N__47458\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47454\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47451\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47449\ : std_logic;
signal \N__47448\ : std_logic;
signal \N__47447\ : std_logic;
signal \N__47446\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47444\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47441\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47438\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47435\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47432\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47424\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47421\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47417\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47091\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47088\ : std_logic;
signal \N__47087\ : std_logic;
signal \N__47086\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47083\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47080\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47077\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47067\ : std_logic;
signal \N__47066\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47063\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47054\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47051\ : std_logic;
signal \N__47050\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47016\ : std_logic;
signal \N__47015\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47010\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47005\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__47002\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46999\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46997\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46994\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46985\ : std_logic;
signal \N__46984\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46982\ : std_logic;
signal \N__46981\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46978\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46973\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46967\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46662\ : std_logic;
signal \N__46659\ : std_logic;
signal \N__46656\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46652\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46650\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46623\ : std_logic;
signal \N__46620\ : std_logic;
signal \N__46613\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46593\ : std_logic;
signal \N__46592\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46568\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46559\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46521\ : std_logic;
signal \N__46512\ : std_logic;
signal \N__46509\ : std_logic;
signal \N__46506\ : std_logic;
signal \N__46503\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46498\ : std_logic;
signal \N__46493\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46481\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46475\ : std_logic;
signal \N__46470\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46466\ : std_logic;
signal \N__46463\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46457\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46449\ : std_logic;
signal \N__46446\ : std_logic;
signal \N__46443\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46434\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46430\ : std_logic;
signal \N__46425\ : std_logic;
signal \N__46420\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46388\ : std_logic;
signal \N__46385\ : std_logic;
signal \N__46382\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46357\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46353\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46345\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46320\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46318\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46312\ : std_logic;
signal \N__46309\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46301\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46295\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46268\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46248\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46230\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46204\ : std_logic;
signal \N__46201\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46182\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46171\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46147\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46104\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46076\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46023\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46004\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45963\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45957\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45946\ : std_logic;
signal \N__45943\ : std_logic;
signal \N__45940\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45922\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45894\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45885\ : std_logic;
signal \N__45882\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45864\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45855\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45851\ : std_logic;
signal \N__45848\ : std_logic;
signal \N__45845\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45813\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45783\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45778\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45761\ : std_logic;
signal \N__45758\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45737\ : std_logic;
signal \N__45734\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45720\ : std_logic;
signal \N__45717\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45687\ : std_logic;
signal \N__45684\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45666\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45654\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45637\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45612\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45597\ : std_logic;
signal \N__45596\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45586\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45566\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45557\ : std_logic;
signal \N__45554\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45542\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45533\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45527\ : std_logic;
signal \N__45524\ : std_logic;
signal \N__45521\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45517\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45480\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45475\ : std_logic;
signal \N__45472\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45424\ : std_logic;
signal \N__45421\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45398\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45378\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45374\ : std_logic;
signal \N__45371\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45369\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45355\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45345\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45340\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45323\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45316\ : std_logic;
signal \N__45313\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45284\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45275\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45262\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45238\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45223\ : std_logic;
signal \N__45220\ : std_logic;
signal \N__45215\ : std_logic;
signal \N__45210\ : std_logic;
signal \N__45207\ : std_logic;
signal \N__45204\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45193\ : std_logic;
signal \N__45188\ : std_logic;
signal \N__45185\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45165\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45158\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45141\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45134\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45122\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45116\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45093\ : std_logic;
signal \N__45092\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45037\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45024\ : std_logic;
signal \N__45021\ : std_logic;
signal \N__45018\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45012\ : std_logic;
signal \N__45011\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44996\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44990\ : std_logic;
signal \N__44987\ : std_logic;
signal \N__44984\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44977\ : std_logic;
signal \N__44976\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44962\ : std_logic;
signal \N__44957\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44940\ : std_logic;
signal \N__44937\ : std_logic;
signal \N__44934\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44921\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44885\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44881\ : std_logic;
signal \N__44878\ : std_logic;
signal \N__44875\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44859\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44842\ : std_logic;
signal \N__44839\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44830\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44808\ : std_logic;
signal \N__44807\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44805\ : std_logic;
signal \N__44802\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44784\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44774\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44768\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44743\ : std_logic;
signal \N__44740\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44727\ : std_logic;
signal \N__44724\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44716\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44701\ : std_logic;
signal \N__44698\ : std_logic;
signal \N__44695\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44673\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44652\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44642\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44638\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44622\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44607\ : std_logic;
signal \N__44604\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44570\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44558\ : std_logic;
signal \N__44555\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44544\ : std_logic;
signal \N__44543\ : std_logic;
signal \N__44540\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44528\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44516\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44498\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44495\ : std_logic;
signal \N__44494\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44492\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44489\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44485\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44483\ : std_logic;
signal \N__44482\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44480\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44475\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44471\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44420\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44393\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44357\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44352\ : std_logic;
signal \N__44349\ : std_logic;
signal \N__44346\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44308\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44297\ : std_logic;
signal \N__44296\ : std_logic;
signal \N__44293\ : std_logic;
signal \N__44290\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44286\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44278\ : std_logic;
signal \N__44275\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44269\ : std_logic;
signal \N__44266\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44248\ : std_logic;
signal \N__44245\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44234\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44230\ : std_logic;
signal \N__44227\ : std_logic;
signal \N__44224\ : std_logic;
signal \N__44221\ : std_logic;
signal \N__44218\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44200\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44159\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44144\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44129\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44120\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44114\ : std_logic;
signal \N__44111\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44100\ : std_logic;
signal \N__44097\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44072\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44057\ : std_logic;
signal \N__44054\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44044\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44036\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44015\ : std_logic;
signal \N__44014\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43995\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43978\ : std_logic;
signal \N__43975\ : std_logic;
signal \N__43972\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43929\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43919\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43907\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43895\ : std_logic;
signal \N__43892\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43860\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43856\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43850\ : std_logic;
signal \N__43845\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43835\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43827\ : std_logic;
signal \N__43826\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43815\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43811\ : std_logic;
signal \N__43808\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43800\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43766\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43762\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43751\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43718\ : std_logic;
signal \N__43713\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43702\ : std_logic;
signal \N__43699\ : std_logic;
signal \N__43696\ : std_logic;
signal \N__43693\ : std_logic;
signal \N__43690\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43672\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43663\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43653\ : std_logic;
signal \N__43650\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43640\ : std_logic;
signal \N__43639\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43608\ : std_logic;
signal \N__43607\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43601\ : std_logic;
signal \N__43598\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43590\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43568\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43554\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43547\ : std_logic;
signal \N__43544\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43509\ : std_logic;
signal \N__43506\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43476\ : std_logic;
signal \N__43473\ : std_logic;
signal \N__43472\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43446\ : std_logic;
signal \N__43443\ : std_logic;
signal \N__43440\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43427\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43416\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43408\ : std_logic;
signal \N__43405\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43391\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43373\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43369\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43353\ : std_logic;
signal \N__43352\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43346\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43334\ : std_logic;
signal \N__43331\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43323\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43312\ : std_logic;
signal \N__43307\ : std_logic;
signal \N__43304\ : std_logic;
signal \N__43303\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43270\ : std_logic;
signal \N__43267\ : std_logic;
signal \N__43264\ : std_logic;
signal \N__43261\ : std_logic;
signal \N__43258\ : std_logic;
signal \N__43255\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43231\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43226\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43203\ : std_logic;
signal \N__43200\ : std_logic;
signal \N__43197\ : std_logic;
signal \N__43194\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43166\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43156\ : std_logic;
signal \N__43153\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43133\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43126\ : std_logic;
signal \N__43123\ : std_logic;
signal \N__43120\ : std_logic;
signal \N__43115\ : std_logic;
signal \N__43114\ : std_logic;
signal \N__43111\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43087\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43078\ : std_logic;
signal \N__43075\ : std_logic;
signal \N__43070\ : std_logic;
signal \N__43069\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43063\ : std_logic;
signal \N__43060\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43046\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43042\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43021\ : std_logic;
signal \N__43018\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42981\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42977\ : std_logic;
signal \N__42974\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42932\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42925\ : std_logic;
signal \N__42922\ : std_logic;
signal \N__42917\ : std_logic;
signal \N__42914\ : std_logic;
signal \N__42913\ : std_logic;
signal \N__42910\ : std_logic;
signal \N__42907\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42894\ : std_logic;
signal \N__42893\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42883\ : std_logic;
signal \N__42880\ : std_logic;
signal \N__42875\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42869\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42851\ : std_logic;
signal \N__42848\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42842\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42832\ : std_logic;
signal \N__42829\ : std_logic;
signal \N__42826\ : std_logic;
signal \N__42821\ : std_logic;
signal \N__42820\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42796\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42781\ : std_logic;
signal \N__42778\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42769\ : std_logic;
signal \N__42766\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42756\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42749\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42736\ : std_logic;
signal \N__42733\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42722\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42709\ : std_logic;
signal \N__42706\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42685\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42672\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42652\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42614\ : std_logic;
signal \N__42613\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42585\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42576\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42568\ : std_logic;
signal \N__42565\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42557\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42546\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42513\ : std_logic;
signal \N__42510\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42504\ : std_logic;
signal \N__42501\ : std_logic;
signal \N__42498\ : std_logic;
signal \N__42495\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42488\ : std_logic;
signal \N__42487\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42469\ : std_logic;
signal \N__42466\ : std_logic;
signal \N__42463\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42449\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42427\ : std_logic;
signal \N__42424\ : std_logic;
signal \N__42421\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42411\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42407\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42400\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42374\ : std_logic;
signal \N__42371\ : std_logic;
signal \N__42368\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42359\ : std_logic;
signal \N__42356\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42296\ : std_logic;
signal \N__42293\ : std_logic;
signal \N__42290\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42284\ : std_logic;
signal \N__42283\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42271\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42255\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42246\ : std_logic;
signal \N__42243\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42231\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42206\ : std_logic;
signal \N__42203\ : std_logic;
signal \N__42200\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42190\ : std_logic;
signal \N__42187\ : std_logic;
signal \N__42184\ : std_logic;
signal \N__42181\ : std_logic;
signal \N__42174\ : std_logic;
signal \N__42171\ : std_logic;
signal \N__42168\ : std_logic;
signal \N__42165\ : std_logic;
signal \N__42162\ : std_logic;
signal \N__42159\ : std_logic;
signal \N__42156\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42122\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42115\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42112\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42109\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42107\ : std_logic;
signal \N__42106\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42104\ : std_logic;
signal \N__42103\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42101\ : std_logic;
signal \N__42100\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42098\ : std_logic;
signal \N__42097\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42094\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42092\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42070\ : std_logic;
signal \N__42061\ : std_logic;
signal \N__42052\ : std_logic;
signal \N__42043\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41997\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41984\ : std_logic;
signal \N__41981\ : std_logic;
signal \N__41978\ : std_logic;
signal \N__41975\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41951\ : std_logic;
signal \N__41948\ : std_logic;
signal \N__41945\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41941\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41927\ : std_logic;
signal \N__41924\ : std_logic;
signal \N__41921\ : std_logic;
signal \N__41918\ : std_logic;
signal \N__41915\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41834\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41798\ : std_logic;
signal \N__41795\ : std_logic;
signal \N__41792\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41756\ : std_logic;
signal \N__41755\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41712\ : std_logic;
signal \N__41709\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41707\ : std_logic;
signal \N__41704\ : std_logic;
signal \N__41699\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41693\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41667\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41657\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41637\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41632\ : std_logic;
signal \N__41627\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41621\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41607\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41573\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41543\ : std_logic;
signal \N__41542\ : std_logic;
signal \N__41537\ : std_logic;
signal \N__41534\ : std_logic;
signal \N__41531\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41504\ : std_logic;
signal \N__41499\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41495\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41489\ : std_logic;
signal \N__41486\ : std_logic;
signal \N__41483\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41459\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41444\ : std_logic;
signal \N__41441\ : std_logic;
signal \N__41438\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41423\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41412\ : std_logic;
signal \N__41409\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41361\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41346\ : std_logic;
signal \N__41345\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41334\ : std_logic;
signal \N__41331\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41290\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41282\ : std_logic;
signal \N__41281\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41258\ : std_logic;
signal \N__41255\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41232\ : std_logic;
signal \N__41229\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41220\ : std_logic;
signal \N__41217\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41192\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41187\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41184\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41174\ : std_logic;
signal \N__41173\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41171\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41168\ : std_logic;
signal \N__41167\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41162\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41159\ : std_logic;
signal \N__41156\ : std_logic;
signal \N__41147\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41137\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41128\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41111\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41105\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41096\ : std_logic;
signal \N__41095\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41092\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41063\ : std_logic;
signal \N__41060\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41045\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41018\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40999\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40995\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40992\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40990\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40964\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40956\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40953\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40950\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40941\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40933\ : std_logic;
signal \N__40930\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40886\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40873\ : std_logic;
signal \N__40870\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40837\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40821\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40755\ : std_logic;
signal \N__40752\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40716\ : std_logic;
signal \N__40715\ : std_logic;
signal \N__40712\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40692\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40662\ : std_logic;
signal \N__40659\ : std_logic;
signal \N__40658\ : std_logic;
signal \N__40655\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40643\ : std_logic;
signal \N__40640\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40628\ : std_logic;
signal \N__40627\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40625\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40613\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40610\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40598\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40595\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40583\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40580\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40565\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40531\ : std_logic;
signal \N__40528\ : std_logic;
signal \N__40519\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40502\ : std_logic;
signal \N__40487\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40484\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40466\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40444\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40442\ : std_logic;
signal \N__40441\ : std_logic;
signal \N__40438\ : std_logic;
signal \N__40435\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40423\ : std_logic;
signal \N__40420\ : std_logic;
signal \N__40417\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40393\ : std_logic;
signal \N__40388\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40363\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40351\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40319\ : std_logic;
signal \N__40312\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40292\ : std_logic;
signal \N__40291\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40270\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40268\ : std_logic;
signal \N__40267\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40265\ : std_logic;
signal \N__40264\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40262\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40246\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40238\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40235\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40232\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40228\ : std_logic;
signal \N__40225\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40208\ : std_logic;
signal \N__40205\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40202\ : std_logic;
signal \N__40201\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40199\ : std_logic;
signal \N__40198\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40196\ : std_logic;
signal \N__40195\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40187\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40175\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40157\ : std_logic;
signal \N__40154\ : std_logic;
signal \N__40151\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40145\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40136\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40133\ : std_logic;
signal \N__40130\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40127\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40121\ : std_logic;
signal \N__40120\ : std_logic;
signal \N__40115\ : std_logic;
signal \N__40114\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40106\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40073\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40052\ : std_logic;
signal \N__40043\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40035\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40029\ : std_logic;
signal \N__40026\ : std_logic;
signal \N__40025\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40016\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40007\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39992\ : std_logic;
signal \N__39989\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39974\ : std_logic;
signal \N__39973\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39970\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39965\ : std_logic;
signal \N__39962\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39956\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39901\ : std_logic;
signal \N__39884\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39808\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39803\ : std_logic;
signal \N__39802\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39785\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39713\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39651\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39630\ : std_logic;
signal \N__39627\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39609\ : std_logic;
signal \N__39606\ : std_logic;
signal \N__39603\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39599\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39583\ : std_logic;
signal \N__39580\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39575\ : std_logic;
signal \N__39572\ : std_logic;
signal \N__39569\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39531\ : std_logic;
signal \N__39528\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39510\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39490\ : std_logic;
signal \N__39487\ : std_logic;
signal \N__39484\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39453\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39444\ : std_logic;
signal \N__39441\ : std_logic;
signal \N__39438\ : std_logic;
signal \N__39437\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39271\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39257\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39251\ : std_logic;
signal \N__39248\ : std_logic;
signal \N__39243\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39232\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39224\ : std_logic;
signal \N__39221\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39215\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39203\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39197\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39185\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39179\ : std_logic;
signal \N__39176\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39163\ : std_logic;
signal \N__39158\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39104\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39080\ : std_logic;
signal \N__39077\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39053\ : std_logic;
signal \N__39050\ : std_logic;
signal \N__39045\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39041\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39024\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39017\ : std_logic;
signal \N__39014\ : std_logic;
signal \N__39009\ : std_logic;
signal \N__39006\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38996\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38987\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38978\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38945\ : std_logic;
signal \N__38942\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38933\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38927\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38915\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38819\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38789\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38783\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38775\ : std_logic;
signal \N__38772\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38616\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38592\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38586\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38517\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38511\ : std_logic;
signal \N__38508\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38478\ : std_logic;
signal \N__38475\ : std_logic;
signal \N__38472\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38448\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38438\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38424\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38361\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38331\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38324\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38289\ : std_logic;
signal \N__38286\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38247\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38225\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38204\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38177\ : std_logic;
signal \N__38174\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38167\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38158\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38114\ : std_logic;
signal \N__38111\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38105\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38063\ : std_logic;
signal \N__38060\ : std_logic;
signal \N__38057\ : std_logic;
signal \N__38054\ : std_logic;
signal \N__38051\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38014\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38011\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38006\ : std_logic;
signal \N__38005\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38003\ : std_logic;
signal \N__38002\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37958\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37916\ : std_logic;
signal \N__37915\ : std_logic;
signal \N__37912\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37896\ : std_logic;
signal \N__37893\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37859\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37828\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37822\ : std_logic;
signal \N__37819\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37741\ : std_logic;
signal \N__37738\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37730\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37708\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37681\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37600\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37578\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37573\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37567\ : std_logic;
signal \N__37564\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37544\ : std_logic;
signal \N__37541\ : std_logic;
signal \N__37538\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37495\ : std_logic;
signal \N__37492\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37471\ : std_logic;
signal \N__37468\ : std_logic;
signal \N__37465\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37423\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37373\ : std_logic;
signal \N__37372\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37354\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37196\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37183\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37112\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37015\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36971\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36916\ : std_logic;
signal \N__36913\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36805\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36730\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36684\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36666\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36536\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36488\ : std_logic;
signal \N__36485\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36461\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36424\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36326\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36320\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36258\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36240\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36175\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36169\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36142\ : std_logic;
signal \N__36139\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36005\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35953\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35950\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35936\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35842\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35836\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35747\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35598\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35595\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35592\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35588\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35529\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35521\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35489\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35423\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35393\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34842\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34341\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34205\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34072\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34028\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34007\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33860\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33788\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33542\ : std_logic;
signal \N__33539\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33344\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33007\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32820\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32749\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32713\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32678\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32642\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32628\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32481\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32478\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32449\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32342\ : std_logic;
signal \N__32339\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32243\ : std_logic;
signal \N__32240\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32053\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31994\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31961\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31463\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31331\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31304\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31271\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31127\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31067\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31055\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31047\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31007\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30947\ : std_logic;
signal \N__30944\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30692\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30614\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30356\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30215\ : std_logic;
signal \N__30212\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29907\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29355\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29343\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29067\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29019\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29004\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28836\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28578\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28523\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27446\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27431\ : std_logic;
signal \N__27428\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27094\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27057\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26905\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25923\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25727\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25658\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25436\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24218\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22868\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20553\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \N_38_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_159\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal pwm_duty_input_0 : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal \pwm_generator_inst.un1_duty_inputlt3\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\ : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\ : std_logic;
signal pwm_duty_input_4 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \rgb_drv_RNOZ0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\ : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \bfn_7_28_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_18\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal s4_phy_c : std_logic;
signal \GB_BUFFER_clock_output_0_THRU_CO\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_198_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_199_i\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.N_1288_i\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_10_26_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_10_27_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \bfn_10_28_0_\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal s3_phy_c : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \bfn_11_24_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \bfn_11_25_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_12_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_12_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_12_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \bfn_12_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal s1_phy_c : std_logic;
signal state_3 : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\ : std_logic;
signal \pll_inst.red_c_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal start_stop_c : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal \bfn_13_22_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.state_RNIE87FZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_13_24_0_\ : std_logic;
signal \pwm_generator_inst.un14_counter_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_13_25_0_\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_201_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_14_20_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal state_ns_i_a3_1 : std_logic;
signal \T45_c\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.time_passed_RNIG7JF\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_200_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_df30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \bfn_15_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_15_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.state_RNI9M3OZ0Z_0\ : std_logic;
signal \phase_controller_inst2.start_timer_tr_RNO_0_0\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \T12_c\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_16_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \T01_c\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \T23_c\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_df30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i_g\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_163_i\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal phase_controller_inst1_state_4 : std_logic;
signal \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\ : std_logic;
signal \phase_controller_inst1.state_RNI7NN7Z0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal clock_output_0 : std_logic;
signal red_c_g : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal clock_output_wire : std_logic;
signal \T01_wire\ : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal \T23_wire\ : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal \T12_wire\ : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal \T45_wire\ : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    clock_output <= clock_output_wire;
    T01 <= \T01_wire\;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    T23 <= \T23_wire\;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    T12 <= \T12_wire\;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    T45 <= \T45_wire\;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__23152\&\N__23160\&\N__23151\&\N__23158\&\N__23150\&\N__23157\&\N__23149\&\N__23159\&\N__23146\&\N__23153\&\N__23145\&\N__23154\&\N__23148\&\N__23155\&\N__23147\&\N__23156\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35583\&'0'&\N__35582\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__36015\&\N__36008\&\N__36013\&\N__36007\&\N__36014\&\N__36006\&\N__36016\&\N__36003\&\N__36009\&\N__36002\&\N__36010\&\N__36004\&\N__36011\&\N__36005\&\N__36012\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35663\&\N__35660\&'0'&'0'&'0'&\N__35658\&\N__35662\&\N__35659\&\N__35661\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__36017\&\N__36020\&\N__36018\&\N__36021\&\N__36019\&\N__19758\&\N__19806\&\N__19824\&\N__19785\&\N__20055\&\N__20105\&\N__20078\&\N__19842\&\N__19857\&\N__19875\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35597\&\N__35594\&'0'&'0'&'0'&\N__35592\&\N__35596\&\N__35593\&\N__35595\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__23110\&\N__22875\&\N__22899\&\N__22926\&\N__22953\&\N__23067\&\N__22977\&\N__23004\&\N__23031\&\N__22434\&\N__22466\&\N__22494\&\N__22518\&\N__22539\&\N__24387\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35670\&'0'&\N__35669\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__24459\,
            RESETB => \N__32172\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clock_output_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__35676\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__35581\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__35664\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__35657\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__35607\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__35591\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__35671\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__35668\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__48637\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48639\,
            DIN => \N__48638\,
            DOUT => \N__48637\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48639\,
            PADOUT => \N__48638\,
            PADIN => \N__48637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48628\,
            DIN => \N__48627\,
            DOUT => \N__48626\,
            PACKAGEPIN => clock_output_wire
        );

    \clock_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48628\,
            PADOUT => \N__48627\,
            PADIN => \N__48626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24477\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T01_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48619\,
            DIN => \N__48618\,
            DOUT => \N__48617\,
            PACKAGEPIN => \T01_wire\
        );

    \T01_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48619\,
            PADOUT => \N__48618\,
            PADIN => \N__48617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__39537\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48610\,
            DIN => \N__48609\,
            DOUT => \N__48608\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48610\,
            PADOUT => \N__48609\,
            PADIN => \N__48608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48601\,
            DIN => \N__48600\,
            DOUT => \N__48599\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48601\,
            PADOUT => \N__48600\,
            PADIN => \N__48599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T23_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48592\,
            DIN => \N__48591\,
            DOUT => \N__48590\,
            PACKAGEPIN => \T23_wire\
        );

    \T23_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48592\,
            PADOUT => \N__48591\,
            PADIN => \N__48590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__41892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48583\,
            DIN => \N__48582\,
            DOUT => \N__48581\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48583\,
            PADOUT => \N__48582\,
            PADIN => \N__48581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33489\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48574\,
            DIN => \N__48573\,
            DOUT => \N__48572\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48574\,
            PADOUT => \N__48573\,
            PADIN => \N__48572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48565\,
            DIN => \N__48564\,
            DOUT => \N__48563\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48565\,
            PADOUT => \N__48564\,
            PADIN => \N__48563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T12_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48556\,
            DIN => \N__48555\,
            DOUT => \N__48554\,
            PACKAGEPIN => \T12_wire\
        );

    \T12_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48556\,
            PADOUT => \N__48555\,
            PADIN => \N__48554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__38433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48547\,
            DIN => \N__48546\,
            DOUT => \N__48545\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48547\,
            PADOUT => \N__48546\,
            PADIN => \N__48545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48538\,
            DIN => \N__48537\,
            DOUT => \N__48536\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48538\,
            PADOUT => \N__48537\,
            PADIN => \N__48536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48529\,
            DIN => \N__48528\,
            DOUT => \N__48527\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48529\,
            PADOUT => \N__48528\,
            PADIN => \N__48527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24360\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48520\,
            DIN => \N__48519\,
            DOUT => \N__48518\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48520\,
            PADOUT => \N__48519\,
            PADIN => \N__48518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48511\,
            DIN => \N__48510\,
            DOUT => \N__48509\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48511\,
            PADOUT => \N__48510\,
            PADIN => \N__48509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29403\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \T45_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48502\,
            DIN => \N__48501\,
            DOUT => \N__48500\,
            PACKAGEPIN => \T45_wire\
        );

    \T45_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__48502\,
            PADOUT => \N__48501\,
            PADIN => \N__48500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48493\,
            DIN => \N__48492\,
            DOUT => \N__48491\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48493\,
            PADOUT => \N__48492\,
            PADIN => \N__48491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__48484\,
            DIN => \N__48483\,
            DOUT => \N__48482\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__48484\,
            PADOUT => \N__48483\,
            PADIN => \N__48482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__11559\ : InMux
    port map (
            O => \N__48465\,
            I => \N__48460\
        );

    \I__11558\ : InMux
    port map (
            O => \N__48464\,
            I => \N__48457\
        );

    \I__11557\ : InMux
    port map (
            O => \N__48463\,
            I => \N__48454\
        );

    \I__11556\ : LocalMux
    port map (
            O => \N__48460\,
            I => \N__48449\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__48457\,
            I => \N__48449\
        );

    \I__11554\ : LocalMux
    port map (
            O => \N__48454\,
            I => \N__48445\
        );

    \I__11553\ : Span4Mux_v
    port map (
            O => \N__48449\,
            I => \N__48442\
        );

    \I__11552\ : InMux
    port map (
            O => \N__48448\,
            I => \N__48439\
        );

    \I__11551\ : Span4Mux_v
    port map (
            O => \N__48445\,
            I => \N__48436\
        );

    \I__11550\ : Sp12to4
    port map (
            O => \N__48442\,
            I => \N__48431\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__48439\,
            I => \N__48431\
        );

    \I__11548\ : Odrv4
    port map (
            O => \N__48436\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__11547\ : Odrv12
    port map (
            O => \N__48431\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__11546\ : InMux
    port map (
            O => \N__48426\,
            I => \N__48422\
        );

    \I__11545\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48418\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__48422\,
            I => \N__48415\
        );

    \I__11543\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48412\
        );

    \I__11542\ : LocalMux
    port map (
            O => \N__48418\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__11541\ : Odrv12
    port map (
            O => \N__48415\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__48412\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__11539\ : InMux
    port map (
            O => \N__48405\,
            I => \N__48402\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__48402\,
            I => \N__48397\
        );

    \I__11537\ : InMux
    port map (
            O => \N__48401\,
            I => \N__48394\
        );

    \I__11536\ : InMux
    port map (
            O => \N__48400\,
            I => \N__48391\
        );

    \I__11535\ : Span4Mux_v
    port map (
            O => \N__48397\,
            I => \N__48388\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__48394\,
            I => \N__48385\
        );

    \I__11533\ : LocalMux
    port map (
            O => \N__48391\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__11532\ : Odrv4
    port map (
            O => \N__48388\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__11531\ : Odrv4
    port map (
            O => \N__48385\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__11530\ : InMux
    port map (
            O => \N__48378\,
            I => \N__48373\
        );

    \I__11529\ : InMux
    port map (
            O => \N__48377\,
            I => \N__48370\
        );

    \I__11528\ : InMux
    port map (
            O => \N__48376\,
            I => \N__48367\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48362\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__48370\,
            I => \N__48362\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__48367\,
            I => \N__48359\
        );

    \I__11524\ : Span12Mux_h
    port map (
            O => \N__48362\,
            I => \N__48355\
        );

    \I__11523\ : Span4Mux_h
    port map (
            O => \N__48359\,
            I => \N__48352\
        );

    \I__11522\ : InMux
    port map (
            O => \N__48358\,
            I => \N__48349\
        );

    \I__11521\ : Odrv12
    port map (
            O => \N__48355\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__11520\ : Odrv4
    port map (
            O => \N__48352\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__48349\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__11518\ : InMux
    port map (
            O => \N__48342\,
            I => \N__48315\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48341\,
            I => \N__48315\
        );

    \I__11516\ : InMux
    port map (
            O => \N__48340\,
            I => \N__48315\
        );

    \I__11515\ : CascadeMux
    port map (
            O => \N__48339\,
            I => \N__48311\
        );

    \I__11514\ : InMux
    port map (
            O => \N__48338\,
            I => \N__48302\
        );

    \I__11513\ : InMux
    port map (
            O => \N__48337\,
            I => \N__48279\
        );

    \I__11512\ : InMux
    port map (
            O => \N__48336\,
            I => \N__48279\
        );

    \I__11511\ : InMux
    port map (
            O => \N__48335\,
            I => \N__48272\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48334\,
            I => \N__48272\
        );

    \I__11509\ : InMux
    port map (
            O => \N__48333\,
            I => \N__48272\
        );

    \I__11508\ : InMux
    port map (
            O => \N__48332\,
            I => \N__48269\
        );

    \I__11507\ : InMux
    port map (
            O => \N__48331\,
            I => \N__48234\
        );

    \I__11506\ : InMux
    port map (
            O => \N__48330\,
            I => \N__48234\
        );

    \I__11505\ : InMux
    port map (
            O => \N__48329\,
            I => \N__48234\
        );

    \I__11504\ : InMux
    port map (
            O => \N__48328\,
            I => \N__48234\
        );

    \I__11503\ : InMux
    port map (
            O => \N__48327\,
            I => \N__48234\
        );

    \I__11502\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48234\
        );

    \I__11501\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48231\
        );

    \I__11500\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48220\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48323\,
            I => \N__48220\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48322\,
            I => \N__48217\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__48315\,
            I => \N__48214\
        );

    \I__11496\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48201\
        );

    \I__11495\ : InMux
    port map (
            O => \N__48311\,
            I => \N__48201\
        );

    \I__11494\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48201\
        );

    \I__11493\ : InMux
    port map (
            O => \N__48309\,
            I => \N__48201\
        );

    \I__11492\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48201\
        );

    \I__11491\ : InMux
    port map (
            O => \N__48307\,
            I => \N__48201\
        );

    \I__11490\ : InMux
    port map (
            O => \N__48306\,
            I => \N__48196\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48305\,
            I => \N__48196\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__48302\,
            I => \N__48193\
        );

    \I__11487\ : InMux
    port map (
            O => \N__48301\,
            I => \N__48173\
        );

    \I__11486\ : InMux
    port map (
            O => \N__48300\,
            I => \N__48173\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48299\,
            I => \N__48173\
        );

    \I__11484\ : InMux
    port map (
            O => \N__48298\,
            I => \N__48173\
        );

    \I__11483\ : InMux
    port map (
            O => \N__48297\,
            I => \N__48173\
        );

    \I__11482\ : InMux
    port map (
            O => \N__48296\,
            I => \N__48166\
        );

    \I__11481\ : InMux
    port map (
            O => \N__48295\,
            I => \N__48166\
        );

    \I__11480\ : InMux
    port map (
            O => \N__48294\,
            I => \N__48166\
        );

    \I__11479\ : InMux
    port map (
            O => \N__48293\,
            I => \N__48163\
        );

    \I__11478\ : InMux
    port map (
            O => \N__48292\,
            I => \N__48152\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48291\,
            I => \N__48152\
        );

    \I__11476\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48152\
        );

    \I__11475\ : InMux
    port map (
            O => \N__48289\,
            I => \N__48152\
        );

    \I__11474\ : InMux
    port map (
            O => \N__48288\,
            I => \N__48152\
        );

    \I__11473\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48143\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48143\
        );

    \I__11471\ : InMux
    port map (
            O => \N__48285\,
            I => \N__48143\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48143\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__48279\,
            I => \N__48138\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__48272\,
            I => \N__48138\
        );

    \I__11467\ : LocalMux
    port map (
            O => \N__48269\,
            I => \N__48135\
        );

    \I__11466\ : InMux
    port map (
            O => \N__48268\,
            I => \N__48132\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48121\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48266\,
            I => \N__48121\
        );

    \I__11463\ : InMux
    port map (
            O => \N__48265\,
            I => \N__48121\
        );

    \I__11462\ : InMux
    port map (
            O => \N__48264\,
            I => \N__48121\
        );

    \I__11461\ : InMux
    port map (
            O => \N__48263\,
            I => \N__48121\
        );

    \I__11460\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48115\
        );

    \I__11459\ : InMux
    port map (
            O => \N__48261\,
            I => \N__48106\
        );

    \I__11458\ : InMux
    port map (
            O => \N__48260\,
            I => \N__48106\
        );

    \I__11457\ : InMux
    port map (
            O => \N__48259\,
            I => \N__48106\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48258\,
            I => \N__48106\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48257\,
            I => \N__48101\
        );

    \I__11454\ : InMux
    port map (
            O => \N__48256\,
            I => \N__48101\
        );

    \I__11453\ : InMux
    port map (
            O => \N__48255\,
            I => \N__48092\
        );

    \I__11452\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48092\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48253\,
            I => \N__48092\
        );

    \I__11450\ : InMux
    port map (
            O => \N__48252\,
            I => \N__48092\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48251\,
            I => \N__48081\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48250\,
            I => \N__48081\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48249\,
            I => \N__48081\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48248\,
            I => \N__48081\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48247\,
            I => \N__48081\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__48234\,
            I => \N__48078\
        );

    \I__11443\ : LocalMux
    port map (
            O => \N__48231\,
            I => \N__48075\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48230\,
            I => \N__48060\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48229\,
            I => \N__48060\
        );

    \I__11440\ : InMux
    port map (
            O => \N__48228\,
            I => \N__48060\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48060\
        );

    \I__11438\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48060\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48225\,
            I => \N__48060\
        );

    \I__11436\ : LocalMux
    port map (
            O => \N__48220\,
            I => \N__48057\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48217\,
            I => \N__48050\
        );

    \I__11434\ : Span4Mux_h
    port map (
            O => \N__48214\,
            I => \N__48050\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__48201\,
            I => \N__48050\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__48196\,
            I => \N__48045\
        );

    \I__11431\ : Span4Mux_v
    port map (
            O => \N__48193\,
            I => \N__48045\
        );

    \I__11430\ : InMux
    port map (
            O => \N__48192\,
            I => \N__48034\
        );

    \I__11429\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48034\
        );

    \I__11428\ : InMux
    port map (
            O => \N__48190\,
            I => \N__48034\
        );

    \I__11427\ : InMux
    port map (
            O => \N__48189\,
            I => \N__48031\
        );

    \I__11426\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48026\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48026\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48019\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48019\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48184\,
            I => \N__48019\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__48173\,
            I => \N__48014\
        );

    \I__11420\ : LocalMux
    port map (
            O => \N__48166\,
            I => \N__48014\
        );

    \I__11419\ : LocalMux
    port map (
            O => \N__48163\,
            I => \N__48011\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__48152\,
            I => \N__48004\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48143\,
            I => \N__48004\
        );

    \I__11416\ : Span4Mux_v
    port map (
            O => \N__48138\,
            I => \N__48004\
        );

    \I__11415\ : Span4Mux_h
    port map (
            O => \N__48135\,
            I => \N__47999\
        );

    \I__11414\ : LocalMux
    port map (
            O => \N__48132\,
            I => \N__47999\
        );

    \I__11413\ : LocalMux
    port map (
            O => \N__48121\,
            I => \N__47996\
        );

    \I__11412\ : InMux
    port map (
            O => \N__48120\,
            I => \N__47993\
        );

    \I__11411\ : InMux
    port map (
            O => \N__48119\,
            I => \N__47988\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48118\,
            I => \N__47988\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__48115\,
            I => \N__47985\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__48106\,
            I => \N__47978\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__47978\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48092\,
            I => \N__47978\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__47971\
        );

    \I__11404\ : Span4Mux_v
    port map (
            O => \N__48078\,
            I => \N__47971\
        );

    \I__11403\ : Span4Mux_v
    port map (
            O => \N__48075\,
            I => \N__47971\
        );

    \I__11402\ : InMux
    port map (
            O => \N__48074\,
            I => \N__47966\
        );

    \I__11401\ : InMux
    port map (
            O => \N__48073\,
            I => \N__47966\
        );

    \I__11400\ : LocalMux
    port map (
            O => \N__48060\,
            I => \N__47957\
        );

    \I__11399\ : Span4Mux_v
    port map (
            O => \N__48057\,
            I => \N__47957\
        );

    \I__11398\ : Span4Mux_v
    port map (
            O => \N__48050\,
            I => \N__47957\
        );

    \I__11397\ : Span4Mux_v
    port map (
            O => \N__48045\,
            I => \N__47957\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48044\,
            I => \N__47954\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48043\,
            I => \N__47947\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48042\,
            I => \N__47947\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48041\,
            I => \N__47947\
        );

    \I__11392\ : LocalMux
    port map (
            O => \N__48034\,
            I => \N__47944\
        );

    \I__11391\ : LocalMux
    port map (
            O => \N__48031\,
            I => \N__47939\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__48026\,
            I => \N__47939\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48019\,
            I => \N__47928\
        );

    \I__11388\ : Span4Mux_v
    port map (
            O => \N__48014\,
            I => \N__47928\
        );

    \I__11387\ : Span4Mux_h
    port map (
            O => \N__48011\,
            I => \N__47928\
        );

    \I__11386\ : Span4Mux_h
    port map (
            O => \N__48004\,
            I => \N__47928\
        );

    \I__11385\ : Span4Mux_h
    port map (
            O => \N__47999\,
            I => \N__47928\
        );

    \I__11384\ : Span12Mux_h
    port map (
            O => \N__47996\,
            I => \N__47925\
        );

    \I__11383\ : LocalMux
    port map (
            O => \N__47993\,
            I => \N__47914\
        );

    \I__11382\ : LocalMux
    port map (
            O => \N__47988\,
            I => \N__47914\
        );

    \I__11381\ : Span4Mux_h
    port map (
            O => \N__47985\,
            I => \N__47914\
        );

    \I__11380\ : Span4Mux_v
    port map (
            O => \N__47978\,
            I => \N__47914\
        );

    \I__11379\ : Span4Mux_h
    port map (
            O => \N__47971\,
            I => \N__47914\
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__47966\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11377\ : Odrv4
    port map (
            O => \N__47957\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11376\ : LocalMux
    port map (
            O => \N__47954\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11375\ : LocalMux
    port map (
            O => \N__47947\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11374\ : Odrv4
    port map (
            O => \N__47944\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11373\ : Odrv4
    port map (
            O => \N__47939\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11372\ : Odrv4
    port map (
            O => \N__47928\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11371\ : Odrv12
    port map (
            O => \N__47925\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11370\ : Odrv4
    port map (
            O => \N__47914\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__11369\ : CascadeMux
    port map (
            O => \N__47895\,
            I => \N__47892\
        );

    \I__11368\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47886\
        );

    \I__11367\ : InMux
    port map (
            O => \N__47891\,
            I => \N__47886\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__47886\,
            I => \N__47883\
        );

    \I__11365\ : Span4Mux_h
    port map (
            O => \N__47883\,
            I => \N__47880\
        );

    \I__11364\ : Odrv4
    port map (
            O => \N__47880\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__11363\ : CEMux
    port map (
            O => \N__47877\,
            I => \N__47870\
        );

    \I__11362\ : CEMux
    port map (
            O => \N__47876\,
            I => \N__47866\
        );

    \I__11361\ : CEMux
    port map (
            O => \N__47875\,
            I => \N__47863\
        );

    \I__11360\ : InMux
    port map (
            O => \N__47874\,
            I => \N__47858\
        );

    \I__11359\ : CEMux
    port map (
            O => \N__47873\,
            I => \N__47855\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__47870\,
            I => \N__47852\
        );

    \I__11357\ : CEMux
    port map (
            O => \N__47869\,
            I => \N__47844\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__47866\,
            I => \N__47816\
        );

    \I__11355\ : LocalMux
    port map (
            O => \N__47863\,
            I => \N__47812\
        );

    \I__11354\ : CEMux
    port map (
            O => \N__47862\,
            I => \N__47808\
        );

    \I__11353\ : CEMux
    port map (
            O => \N__47861\,
            I => \N__47805\
        );

    \I__11352\ : LocalMux
    port map (
            O => \N__47858\,
            I => \N__47802\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__47855\,
            I => \N__47799\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__47852\,
            I => \N__47796\
        );

    \I__11349\ : CEMux
    port map (
            O => \N__47851\,
            I => \N__47793\
        );

    \I__11348\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47784\
        );

    \I__11347\ : InMux
    port map (
            O => \N__47849\,
            I => \N__47784\
        );

    \I__11346\ : InMux
    port map (
            O => \N__47848\,
            I => \N__47784\
        );

    \I__11345\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47784\
        );

    \I__11344\ : LocalMux
    port map (
            O => \N__47844\,
            I => \N__47781\
        );

    \I__11343\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47770\
        );

    \I__11342\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47770\
        );

    \I__11341\ : InMux
    port map (
            O => \N__47841\,
            I => \N__47770\
        );

    \I__11340\ : InMux
    port map (
            O => \N__47840\,
            I => \N__47761\
        );

    \I__11339\ : InMux
    port map (
            O => \N__47839\,
            I => \N__47761\
        );

    \I__11338\ : InMux
    port map (
            O => \N__47838\,
            I => \N__47761\
        );

    \I__11337\ : InMux
    port map (
            O => \N__47837\,
            I => \N__47761\
        );

    \I__11336\ : InMux
    port map (
            O => \N__47836\,
            I => \N__47752\
        );

    \I__11335\ : InMux
    port map (
            O => \N__47835\,
            I => \N__47752\
        );

    \I__11334\ : InMux
    port map (
            O => \N__47834\,
            I => \N__47752\
        );

    \I__11333\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47752\
        );

    \I__11332\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47743\
        );

    \I__11331\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47743\
        );

    \I__11330\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47743\
        );

    \I__11329\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47743\
        );

    \I__11328\ : InMux
    port map (
            O => \N__47828\,
            I => \N__47736\
        );

    \I__11327\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47736\
        );

    \I__11326\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47736\
        );

    \I__11325\ : CEMux
    port map (
            O => \N__47825\,
            I => \N__47732\
        );

    \I__11324\ : CEMux
    port map (
            O => \N__47824\,
            I => \N__47729\
        );

    \I__11323\ : CEMux
    port map (
            O => \N__47823\,
            I => \N__47726\
        );

    \I__11322\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47717\
        );

    \I__11321\ : InMux
    port map (
            O => \N__47821\,
            I => \N__47717\
        );

    \I__11320\ : InMux
    port map (
            O => \N__47820\,
            I => \N__47717\
        );

    \I__11319\ : InMux
    port map (
            O => \N__47819\,
            I => \N__47717\
        );

    \I__11318\ : Span4Mux_v
    port map (
            O => \N__47816\,
            I => \N__47714\
        );

    \I__11317\ : CEMux
    port map (
            O => \N__47815\,
            I => \N__47711\
        );

    \I__11316\ : Span4Mux_v
    port map (
            O => \N__47812\,
            I => \N__47708\
        );

    \I__11315\ : CEMux
    port map (
            O => \N__47811\,
            I => \N__47705\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__47808\,
            I => \N__47702\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__47805\,
            I => \N__47699\
        );

    \I__11312\ : Span4Mux_v
    port map (
            O => \N__47802\,
            I => \N__47696\
        );

    \I__11311\ : Span4Mux_h
    port map (
            O => \N__47799\,
            I => \N__47685\
        );

    \I__11310\ : Span4Mux_h
    port map (
            O => \N__47796\,
            I => \N__47685\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__47793\,
            I => \N__47685\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__47784\,
            I => \N__47685\
        );

    \I__11307\ : Span4Mux_v
    port map (
            O => \N__47781\,
            I => \N__47685\
        );

    \I__11306\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47676\
        );

    \I__11305\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47676\
        );

    \I__11304\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47676\
        );

    \I__11303\ : InMux
    port map (
            O => \N__47777\,
            I => \N__47676\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__47770\,
            I => \N__47671\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__47761\,
            I => \N__47671\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__47752\,
            I => \N__47664\
        );

    \I__11299\ : LocalMux
    port map (
            O => \N__47743\,
            I => \N__47664\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__47736\,
            I => \N__47664\
        );

    \I__11297\ : CEMux
    port map (
            O => \N__47735\,
            I => \N__47661\
        );

    \I__11296\ : LocalMux
    port map (
            O => \N__47732\,
            I => \N__47656\
        );

    \I__11295\ : LocalMux
    port map (
            O => \N__47729\,
            I => \N__47656\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__47726\,
            I => \N__47653\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__47717\,
            I => \N__47648\
        );

    \I__11292\ : Span4Mux_h
    port map (
            O => \N__47714\,
            I => \N__47648\
        );

    \I__11291\ : LocalMux
    port map (
            O => \N__47711\,
            I => \N__47645\
        );

    \I__11290\ : Span4Mux_h
    port map (
            O => \N__47708\,
            I => \N__47640\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__47705\,
            I => \N__47640\
        );

    \I__11288\ : Span4Mux_v
    port map (
            O => \N__47702\,
            I => \N__47635\
        );

    \I__11287\ : Span4Mux_h
    port map (
            O => \N__47699\,
            I => \N__47635\
        );

    \I__11286\ : Span4Mux_h
    port map (
            O => \N__47696\,
            I => \N__47632\
        );

    \I__11285\ : Span4Mux_v
    port map (
            O => \N__47685\,
            I => \N__47623\
        );

    \I__11284\ : LocalMux
    port map (
            O => \N__47676\,
            I => \N__47623\
        );

    \I__11283\ : Span4Mux_v
    port map (
            O => \N__47671\,
            I => \N__47623\
        );

    \I__11282\ : Span4Mux_v
    port map (
            O => \N__47664\,
            I => \N__47623\
        );

    \I__11281\ : LocalMux
    port map (
            O => \N__47661\,
            I => \N__47618\
        );

    \I__11280\ : Span12Mux_h
    port map (
            O => \N__47656\,
            I => \N__47618\
        );

    \I__11279\ : Span4Mux_v
    port map (
            O => \N__47653\,
            I => \N__47613\
        );

    \I__11278\ : Span4Mux_h
    port map (
            O => \N__47648\,
            I => \N__47613\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__47645\,
            I => \N__47610\
        );

    \I__11276\ : Sp12to4
    port map (
            O => \N__47640\,
            I => \N__47607\
        );

    \I__11275\ : Span4Mux_h
    port map (
            O => \N__47635\,
            I => \N__47604\
        );

    \I__11274\ : Span4Mux_h
    port map (
            O => \N__47632\,
            I => \N__47601\
        );

    \I__11273\ : Span4Mux_h
    port map (
            O => \N__47623\,
            I => \N__47598\
        );

    \I__11272\ : Odrv12
    port map (
            O => \N__47618\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11271\ : Odrv4
    port map (
            O => \N__47613\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11270\ : Odrv4
    port map (
            O => \N__47610\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11269\ : Odrv12
    port map (
            O => \N__47607\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11268\ : Odrv4
    port map (
            O => \N__47604\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11267\ : Odrv4
    port map (
            O => \N__47601\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11266\ : Odrv4
    port map (
            O => \N__47598\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__11265\ : InMux
    port map (
            O => \N__47583\,
            I => \N__47580\
        );

    \I__11264\ : LocalMux
    port map (
            O => \N__47580\,
            I => \N__47577\
        );

    \I__11263\ : Span4Mux_v
    port map (
            O => \N__47577\,
            I => \N__47573\
        );

    \I__11262\ : InMux
    port map (
            O => \N__47576\,
            I => \N__47570\
        );

    \I__11261\ : Span4Mux_h
    port map (
            O => \N__47573\,
            I => \N__47567\
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__47570\,
            I => \N__47564\
        );

    \I__11259\ : Odrv4
    port map (
            O => \N__47567\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__11258\ : Odrv4
    port map (
            O => \N__47564\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__11257\ : InMux
    port map (
            O => \N__47559\,
            I => \N__47556\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__47556\,
            I => \N__47413\
        );

    \I__11255\ : ClkMux
    port map (
            O => \N__47555\,
            I => \N__47127\
        );

    \I__11254\ : ClkMux
    port map (
            O => \N__47554\,
            I => \N__47127\
        );

    \I__11253\ : ClkMux
    port map (
            O => \N__47553\,
            I => \N__47127\
        );

    \I__11252\ : ClkMux
    port map (
            O => \N__47552\,
            I => \N__47127\
        );

    \I__11251\ : ClkMux
    port map (
            O => \N__47551\,
            I => \N__47127\
        );

    \I__11250\ : ClkMux
    port map (
            O => \N__47550\,
            I => \N__47127\
        );

    \I__11249\ : ClkMux
    port map (
            O => \N__47549\,
            I => \N__47127\
        );

    \I__11248\ : ClkMux
    port map (
            O => \N__47548\,
            I => \N__47127\
        );

    \I__11247\ : ClkMux
    port map (
            O => \N__47547\,
            I => \N__47127\
        );

    \I__11246\ : ClkMux
    port map (
            O => \N__47546\,
            I => \N__47127\
        );

    \I__11245\ : ClkMux
    port map (
            O => \N__47545\,
            I => \N__47127\
        );

    \I__11244\ : ClkMux
    port map (
            O => \N__47544\,
            I => \N__47127\
        );

    \I__11243\ : ClkMux
    port map (
            O => \N__47543\,
            I => \N__47127\
        );

    \I__11242\ : ClkMux
    port map (
            O => \N__47542\,
            I => \N__47127\
        );

    \I__11241\ : ClkMux
    port map (
            O => \N__47541\,
            I => \N__47127\
        );

    \I__11240\ : ClkMux
    port map (
            O => \N__47540\,
            I => \N__47127\
        );

    \I__11239\ : ClkMux
    port map (
            O => \N__47539\,
            I => \N__47127\
        );

    \I__11238\ : ClkMux
    port map (
            O => \N__47538\,
            I => \N__47127\
        );

    \I__11237\ : ClkMux
    port map (
            O => \N__47537\,
            I => \N__47127\
        );

    \I__11236\ : ClkMux
    port map (
            O => \N__47536\,
            I => \N__47127\
        );

    \I__11235\ : ClkMux
    port map (
            O => \N__47535\,
            I => \N__47127\
        );

    \I__11234\ : ClkMux
    port map (
            O => \N__47534\,
            I => \N__47127\
        );

    \I__11233\ : ClkMux
    port map (
            O => \N__47533\,
            I => \N__47127\
        );

    \I__11232\ : ClkMux
    port map (
            O => \N__47532\,
            I => \N__47127\
        );

    \I__11231\ : ClkMux
    port map (
            O => \N__47531\,
            I => \N__47127\
        );

    \I__11230\ : ClkMux
    port map (
            O => \N__47530\,
            I => \N__47127\
        );

    \I__11229\ : ClkMux
    port map (
            O => \N__47529\,
            I => \N__47127\
        );

    \I__11228\ : ClkMux
    port map (
            O => \N__47528\,
            I => \N__47127\
        );

    \I__11227\ : ClkMux
    port map (
            O => \N__47527\,
            I => \N__47127\
        );

    \I__11226\ : ClkMux
    port map (
            O => \N__47526\,
            I => \N__47127\
        );

    \I__11225\ : ClkMux
    port map (
            O => \N__47525\,
            I => \N__47127\
        );

    \I__11224\ : ClkMux
    port map (
            O => \N__47524\,
            I => \N__47127\
        );

    \I__11223\ : ClkMux
    port map (
            O => \N__47523\,
            I => \N__47127\
        );

    \I__11222\ : ClkMux
    port map (
            O => \N__47522\,
            I => \N__47127\
        );

    \I__11221\ : ClkMux
    port map (
            O => \N__47521\,
            I => \N__47127\
        );

    \I__11220\ : ClkMux
    port map (
            O => \N__47520\,
            I => \N__47127\
        );

    \I__11219\ : ClkMux
    port map (
            O => \N__47519\,
            I => \N__47127\
        );

    \I__11218\ : ClkMux
    port map (
            O => \N__47518\,
            I => \N__47127\
        );

    \I__11217\ : ClkMux
    port map (
            O => \N__47517\,
            I => \N__47127\
        );

    \I__11216\ : ClkMux
    port map (
            O => \N__47516\,
            I => \N__47127\
        );

    \I__11215\ : ClkMux
    port map (
            O => \N__47515\,
            I => \N__47127\
        );

    \I__11214\ : ClkMux
    port map (
            O => \N__47514\,
            I => \N__47127\
        );

    \I__11213\ : ClkMux
    port map (
            O => \N__47513\,
            I => \N__47127\
        );

    \I__11212\ : ClkMux
    port map (
            O => \N__47512\,
            I => \N__47127\
        );

    \I__11211\ : ClkMux
    port map (
            O => \N__47511\,
            I => \N__47127\
        );

    \I__11210\ : ClkMux
    port map (
            O => \N__47510\,
            I => \N__47127\
        );

    \I__11209\ : ClkMux
    port map (
            O => \N__47509\,
            I => \N__47127\
        );

    \I__11208\ : ClkMux
    port map (
            O => \N__47508\,
            I => \N__47127\
        );

    \I__11207\ : ClkMux
    port map (
            O => \N__47507\,
            I => \N__47127\
        );

    \I__11206\ : ClkMux
    port map (
            O => \N__47506\,
            I => \N__47127\
        );

    \I__11205\ : ClkMux
    port map (
            O => \N__47505\,
            I => \N__47127\
        );

    \I__11204\ : ClkMux
    port map (
            O => \N__47504\,
            I => \N__47127\
        );

    \I__11203\ : ClkMux
    port map (
            O => \N__47503\,
            I => \N__47127\
        );

    \I__11202\ : ClkMux
    port map (
            O => \N__47502\,
            I => \N__47127\
        );

    \I__11201\ : ClkMux
    port map (
            O => \N__47501\,
            I => \N__47127\
        );

    \I__11200\ : ClkMux
    port map (
            O => \N__47500\,
            I => \N__47127\
        );

    \I__11199\ : ClkMux
    port map (
            O => \N__47499\,
            I => \N__47127\
        );

    \I__11198\ : ClkMux
    port map (
            O => \N__47498\,
            I => \N__47127\
        );

    \I__11197\ : ClkMux
    port map (
            O => \N__47497\,
            I => \N__47127\
        );

    \I__11196\ : ClkMux
    port map (
            O => \N__47496\,
            I => \N__47127\
        );

    \I__11195\ : ClkMux
    port map (
            O => \N__47495\,
            I => \N__47127\
        );

    \I__11194\ : ClkMux
    port map (
            O => \N__47494\,
            I => \N__47127\
        );

    \I__11193\ : ClkMux
    port map (
            O => \N__47493\,
            I => \N__47127\
        );

    \I__11192\ : ClkMux
    port map (
            O => \N__47492\,
            I => \N__47127\
        );

    \I__11191\ : ClkMux
    port map (
            O => \N__47491\,
            I => \N__47127\
        );

    \I__11190\ : ClkMux
    port map (
            O => \N__47490\,
            I => \N__47127\
        );

    \I__11189\ : ClkMux
    port map (
            O => \N__47489\,
            I => \N__47127\
        );

    \I__11188\ : ClkMux
    port map (
            O => \N__47488\,
            I => \N__47127\
        );

    \I__11187\ : ClkMux
    port map (
            O => \N__47487\,
            I => \N__47127\
        );

    \I__11186\ : ClkMux
    port map (
            O => \N__47486\,
            I => \N__47127\
        );

    \I__11185\ : ClkMux
    port map (
            O => \N__47485\,
            I => \N__47127\
        );

    \I__11184\ : ClkMux
    port map (
            O => \N__47484\,
            I => \N__47127\
        );

    \I__11183\ : ClkMux
    port map (
            O => \N__47483\,
            I => \N__47127\
        );

    \I__11182\ : ClkMux
    port map (
            O => \N__47482\,
            I => \N__47127\
        );

    \I__11181\ : ClkMux
    port map (
            O => \N__47481\,
            I => \N__47127\
        );

    \I__11180\ : ClkMux
    port map (
            O => \N__47480\,
            I => \N__47127\
        );

    \I__11179\ : ClkMux
    port map (
            O => \N__47479\,
            I => \N__47127\
        );

    \I__11178\ : ClkMux
    port map (
            O => \N__47478\,
            I => \N__47127\
        );

    \I__11177\ : ClkMux
    port map (
            O => \N__47477\,
            I => \N__47127\
        );

    \I__11176\ : ClkMux
    port map (
            O => \N__47476\,
            I => \N__47127\
        );

    \I__11175\ : ClkMux
    port map (
            O => \N__47475\,
            I => \N__47127\
        );

    \I__11174\ : ClkMux
    port map (
            O => \N__47474\,
            I => \N__47127\
        );

    \I__11173\ : ClkMux
    port map (
            O => \N__47473\,
            I => \N__47127\
        );

    \I__11172\ : ClkMux
    port map (
            O => \N__47472\,
            I => \N__47127\
        );

    \I__11171\ : ClkMux
    port map (
            O => \N__47471\,
            I => \N__47127\
        );

    \I__11170\ : ClkMux
    port map (
            O => \N__47470\,
            I => \N__47127\
        );

    \I__11169\ : ClkMux
    port map (
            O => \N__47469\,
            I => \N__47127\
        );

    \I__11168\ : ClkMux
    port map (
            O => \N__47468\,
            I => \N__47127\
        );

    \I__11167\ : ClkMux
    port map (
            O => \N__47467\,
            I => \N__47127\
        );

    \I__11166\ : ClkMux
    port map (
            O => \N__47466\,
            I => \N__47127\
        );

    \I__11165\ : ClkMux
    port map (
            O => \N__47465\,
            I => \N__47127\
        );

    \I__11164\ : ClkMux
    port map (
            O => \N__47464\,
            I => \N__47127\
        );

    \I__11163\ : ClkMux
    port map (
            O => \N__47463\,
            I => \N__47127\
        );

    \I__11162\ : ClkMux
    port map (
            O => \N__47462\,
            I => \N__47127\
        );

    \I__11161\ : ClkMux
    port map (
            O => \N__47461\,
            I => \N__47127\
        );

    \I__11160\ : ClkMux
    port map (
            O => \N__47460\,
            I => \N__47127\
        );

    \I__11159\ : ClkMux
    port map (
            O => \N__47459\,
            I => \N__47127\
        );

    \I__11158\ : ClkMux
    port map (
            O => \N__47458\,
            I => \N__47127\
        );

    \I__11157\ : ClkMux
    port map (
            O => \N__47457\,
            I => \N__47127\
        );

    \I__11156\ : ClkMux
    port map (
            O => \N__47456\,
            I => \N__47127\
        );

    \I__11155\ : ClkMux
    port map (
            O => \N__47455\,
            I => \N__47127\
        );

    \I__11154\ : ClkMux
    port map (
            O => \N__47454\,
            I => \N__47127\
        );

    \I__11153\ : ClkMux
    port map (
            O => \N__47453\,
            I => \N__47127\
        );

    \I__11152\ : ClkMux
    port map (
            O => \N__47452\,
            I => \N__47127\
        );

    \I__11151\ : ClkMux
    port map (
            O => \N__47451\,
            I => \N__47127\
        );

    \I__11150\ : ClkMux
    port map (
            O => \N__47450\,
            I => \N__47127\
        );

    \I__11149\ : ClkMux
    port map (
            O => \N__47449\,
            I => \N__47127\
        );

    \I__11148\ : ClkMux
    port map (
            O => \N__47448\,
            I => \N__47127\
        );

    \I__11147\ : ClkMux
    port map (
            O => \N__47447\,
            I => \N__47127\
        );

    \I__11146\ : ClkMux
    port map (
            O => \N__47446\,
            I => \N__47127\
        );

    \I__11145\ : ClkMux
    port map (
            O => \N__47445\,
            I => \N__47127\
        );

    \I__11144\ : ClkMux
    port map (
            O => \N__47444\,
            I => \N__47127\
        );

    \I__11143\ : ClkMux
    port map (
            O => \N__47443\,
            I => \N__47127\
        );

    \I__11142\ : ClkMux
    port map (
            O => \N__47442\,
            I => \N__47127\
        );

    \I__11141\ : ClkMux
    port map (
            O => \N__47441\,
            I => \N__47127\
        );

    \I__11140\ : ClkMux
    port map (
            O => \N__47440\,
            I => \N__47127\
        );

    \I__11139\ : ClkMux
    port map (
            O => \N__47439\,
            I => \N__47127\
        );

    \I__11138\ : ClkMux
    port map (
            O => \N__47438\,
            I => \N__47127\
        );

    \I__11137\ : ClkMux
    port map (
            O => \N__47437\,
            I => \N__47127\
        );

    \I__11136\ : ClkMux
    port map (
            O => \N__47436\,
            I => \N__47127\
        );

    \I__11135\ : ClkMux
    port map (
            O => \N__47435\,
            I => \N__47127\
        );

    \I__11134\ : ClkMux
    port map (
            O => \N__47434\,
            I => \N__47127\
        );

    \I__11133\ : ClkMux
    port map (
            O => \N__47433\,
            I => \N__47127\
        );

    \I__11132\ : ClkMux
    port map (
            O => \N__47432\,
            I => \N__47127\
        );

    \I__11131\ : ClkMux
    port map (
            O => \N__47431\,
            I => \N__47127\
        );

    \I__11130\ : ClkMux
    port map (
            O => \N__47430\,
            I => \N__47127\
        );

    \I__11129\ : ClkMux
    port map (
            O => \N__47429\,
            I => \N__47127\
        );

    \I__11128\ : ClkMux
    port map (
            O => \N__47428\,
            I => \N__47127\
        );

    \I__11127\ : ClkMux
    port map (
            O => \N__47427\,
            I => \N__47127\
        );

    \I__11126\ : ClkMux
    port map (
            O => \N__47426\,
            I => \N__47127\
        );

    \I__11125\ : ClkMux
    port map (
            O => \N__47425\,
            I => \N__47127\
        );

    \I__11124\ : ClkMux
    port map (
            O => \N__47424\,
            I => \N__47127\
        );

    \I__11123\ : ClkMux
    port map (
            O => \N__47423\,
            I => \N__47127\
        );

    \I__11122\ : ClkMux
    port map (
            O => \N__47422\,
            I => \N__47127\
        );

    \I__11121\ : ClkMux
    port map (
            O => \N__47421\,
            I => \N__47127\
        );

    \I__11120\ : ClkMux
    port map (
            O => \N__47420\,
            I => \N__47127\
        );

    \I__11119\ : ClkMux
    port map (
            O => \N__47419\,
            I => \N__47127\
        );

    \I__11118\ : ClkMux
    port map (
            O => \N__47418\,
            I => \N__47127\
        );

    \I__11117\ : ClkMux
    port map (
            O => \N__47417\,
            I => \N__47127\
        );

    \I__11116\ : ClkMux
    port map (
            O => \N__47416\,
            I => \N__47127\
        );

    \I__11115\ : Glb2LocalMux
    port map (
            O => \N__47413\,
            I => \N__47127\
        );

    \I__11114\ : ClkMux
    port map (
            O => \N__47412\,
            I => \N__47127\
        );

    \I__11113\ : GlobalMux
    port map (
            O => \N__47127\,
            I => clock_output_0
        );

    \I__11112\ : InMux
    port map (
            O => \N__47124\,
            I => \N__47118\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47123\,
            I => \N__47115\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47122\,
            I => \N__47112\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47109\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__47118\,
            I => \N__47106\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47115\,
            I => \N__47103\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47112\,
            I => \N__47100\
        );

    \I__11105\ : LocalMux
    port map (
            O => \N__47109\,
            I => \N__47095\
        );

    \I__11104\ : Glb2LocalMux
    port map (
            O => \N__47106\,
            I => \N__46662\
        );

    \I__11103\ : Glb2LocalMux
    port map (
            O => \N__47103\,
            I => \N__46662\
        );

    \I__11102\ : Glb2LocalMux
    port map (
            O => \N__47100\,
            I => \N__46662\
        );

    \I__11101\ : SRMux
    port map (
            O => \N__47099\,
            I => \N__46662\
        );

    \I__11100\ : SRMux
    port map (
            O => \N__47098\,
            I => \N__46662\
        );

    \I__11099\ : Glb2LocalMux
    port map (
            O => \N__47095\,
            I => \N__46662\
        );

    \I__11098\ : SRMux
    port map (
            O => \N__47094\,
            I => \N__46662\
        );

    \I__11097\ : SRMux
    port map (
            O => \N__47093\,
            I => \N__46662\
        );

    \I__11096\ : SRMux
    port map (
            O => \N__47092\,
            I => \N__46662\
        );

    \I__11095\ : SRMux
    port map (
            O => \N__47091\,
            I => \N__46662\
        );

    \I__11094\ : SRMux
    port map (
            O => \N__47090\,
            I => \N__46662\
        );

    \I__11093\ : SRMux
    port map (
            O => \N__47089\,
            I => \N__46662\
        );

    \I__11092\ : SRMux
    port map (
            O => \N__47088\,
            I => \N__46662\
        );

    \I__11091\ : SRMux
    port map (
            O => \N__47087\,
            I => \N__46662\
        );

    \I__11090\ : SRMux
    port map (
            O => \N__47086\,
            I => \N__46662\
        );

    \I__11089\ : SRMux
    port map (
            O => \N__47085\,
            I => \N__46662\
        );

    \I__11088\ : SRMux
    port map (
            O => \N__47084\,
            I => \N__46662\
        );

    \I__11087\ : SRMux
    port map (
            O => \N__47083\,
            I => \N__46662\
        );

    \I__11086\ : SRMux
    port map (
            O => \N__47082\,
            I => \N__46662\
        );

    \I__11085\ : SRMux
    port map (
            O => \N__47081\,
            I => \N__46662\
        );

    \I__11084\ : SRMux
    port map (
            O => \N__47080\,
            I => \N__46662\
        );

    \I__11083\ : SRMux
    port map (
            O => \N__47079\,
            I => \N__46662\
        );

    \I__11082\ : SRMux
    port map (
            O => \N__47078\,
            I => \N__46662\
        );

    \I__11081\ : SRMux
    port map (
            O => \N__47077\,
            I => \N__46662\
        );

    \I__11080\ : SRMux
    port map (
            O => \N__47076\,
            I => \N__46662\
        );

    \I__11079\ : SRMux
    port map (
            O => \N__47075\,
            I => \N__46662\
        );

    \I__11078\ : SRMux
    port map (
            O => \N__47074\,
            I => \N__46662\
        );

    \I__11077\ : SRMux
    port map (
            O => \N__47073\,
            I => \N__46662\
        );

    \I__11076\ : SRMux
    port map (
            O => \N__47072\,
            I => \N__46662\
        );

    \I__11075\ : SRMux
    port map (
            O => \N__47071\,
            I => \N__46662\
        );

    \I__11074\ : SRMux
    port map (
            O => \N__47070\,
            I => \N__46662\
        );

    \I__11073\ : SRMux
    port map (
            O => \N__47069\,
            I => \N__46662\
        );

    \I__11072\ : SRMux
    port map (
            O => \N__47068\,
            I => \N__46662\
        );

    \I__11071\ : SRMux
    port map (
            O => \N__47067\,
            I => \N__46662\
        );

    \I__11070\ : SRMux
    port map (
            O => \N__47066\,
            I => \N__46662\
        );

    \I__11069\ : SRMux
    port map (
            O => \N__47065\,
            I => \N__46662\
        );

    \I__11068\ : SRMux
    port map (
            O => \N__47064\,
            I => \N__46662\
        );

    \I__11067\ : SRMux
    port map (
            O => \N__47063\,
            I => \N__46662\
        );

    \I__11066\ : SRMux
    port map (
            O => \N__47062\,
            I => \N__46662\
        );

    \I__11065\ : SRMux
    port map (
            O => \N__47061\,
            I => \N__46662\
        );

    \I__11064\ : SRMux
    port map (
            O => \N__47060\,
            I => \N__46662\
        );

    \I__11063\ : SRMux
    port map (
            O => \N__47059\,
            I => \N__46662\
        );

    \I__11062\ : SRMux
    port map (
            O => \N__47058\,
            I => \N__46662\
        );

    \I__11061\ : SRMux
    port map (
            O => \N__47057\,
            I => \N__46662\
        );

    \I__11060\ : SRMux
    port map (
            O => \N__47056\,
            I => \N__46662\
        );

    \I__11059\ : SRMux
    port map (
            O => \N__47055\,
            I => \N__46662\
        );

    \I__11058\ : SRMux
    port map (
            O => \N__47054\,
            I => \N__46662\
        );

    \I__11057\ : SRMux
    port map (
            O => \N__47053\,
            I => \N__46662\
        );

    \I__11056\ : SRMux
    port map (
            O => \N__47052\,
            I => \N__46662\
        );

    \I__11055\ : SRMux
    port map (
            O => \N__47051\,
            I => \N__46662\
        );

    \I__11054\ : SRMux
    port map (
            O => \N__47050\,
            I => \N__46662\
        );

    \I__11053\ : SRMux
    port map (
            O => \N__47049\,
            I => \N__46662\
        );

    \I__11052\ : SRMux
    port map (
            O => \N__47048\,
            I => \N__46662\
        );

    \I__11051\ : SRMux
    port map (
            O => \N__47047\,
            I => \N__46662\
        );

    \I__11050\ : SRMux
    port map (
            O => \N__47046\,
            I => \N__46662\
        );

    \I__11049\ : SRMux
    port map (
            O => \N__47045\,
            I => \N__46662\
        );

    \I__11048\ : SRMux
    port map (
            O => \N__47044\,
            I => \N__46662\
        );

    \I__11047\ : SRMux
    port map (
            O => \N__47043\,
            I => \N__46662\
        );

    \I__11046\ : SRMux
    port map (
            O => \N__47042\,
            I => \N__46662\
        );

    \I__11045\ : SRMux
    port map (
            O => \N__47041\,
            I => \N__46662\
        );

    \I__11044\ : SRMux
    port map (
            O => \N__47040\,
            I => \N__46662\
        );

    \I__11043\ : SRMux
    port map (
            O => \N__47039\,
            I => \N__46662\
        );

    \I__11042\ : SRMux
    port map (
            O => \N__47038\,
            I => \N__46662\
        );

    \I__11041\ : SRMux
    port map (
            O => \N__47037\,
            I => \N__46662\
        );

    \I__11040\ : SRMux
    port map (
            O => \N__47036\,
            I => \N__46662\
        );

    \I__11039\ : SRMux
    port map (
            O => \N__47035\,
            I => \N__46662\
        );

    \I__11038\ : SRMux
    port map (
            O => \N__47034\,
            I => \N__46662\
        );

    \I__11037\ : SRMux
    port map (
            O => \N__47033\,
            I => \N__46662\
        );

    \I__11036\ : SRMux
    port map (
            O => \N__47032\,
            I => \N__46662\
        );

    \I__11035\ : SRMux
    port map (
            O => \N__47031\,
            I => \N__46662\
        );

    \I__11034\ : SRMux
    port map (
            O => \N__47030\,
            I => \N__46662\
        );

    \I__11033\ : SRMux
    port map (
            O => \N__47029\,
            I => \N__46662\
        );

    \I__11032\ : SRMux
    port map (
            O => \N__47028\,
            I => \N__46662\
        );

    \I__11031\ : SRMux
    port map (
            O => \N__47027\,
            I => \N__46662\
        );

    \I__11030\ : SRMux
    port map (
            O => \N__47026\,
            I => \N__46662\
        );

    \I__11029\ : SRMux
    port map (
            O => \N__47025\,
            I => \N__46662\
        );

    \I__11028\ : SRMux
    port map (
            O => \N__47024\,
            I => \N__46662\
        );

    \I__11027\ : SRMux
    port map (
            O => \N__47023\,
            I => \N__46662\
        );

    \I__11026\ : SRMux
    port map (
            O => \N__47022\,
            I => \N__46662\
        );

    \I__11025\ : SRMux
    port map (
            O => \N__47021\,
            I => \N__46662\
        );

    \I__11024\ : SRMux
    port map (
            O => \N__47020\,
            I => \N__46662\
        );

    \I__11023\ : SRMux
    port map (
            O => \N__47019\,
            I => \N__46662\
        );

    \I__11022\ : SRMux
    port map (
            O => \N__47018\,
            I => \N__46662\
        );

    \I__11021\ : SRMux
    port map (
            O => \N__47017\,
            I => \N__46662\
        );

    \I__11020\ : SRMux
    port map (
            O => \N__47016\,
            I => \N__46662\
        );

    \I__11019\ : SRMux
    port map (
            O => \N__47015\,
            I => \N__46662\
        );

    \I__11018\ : SRMux
    port map (
            O => \N__47014\,
            I => \N__46662\
        );

    \I__11017\ : SRMux
    port map (
            O => \N__47013\,
            I => \N__46662\
        );

    \I__11016\ : SRMux
    port map (
            O => \N__47012\,
            I => \N__46662\
        );

    \I__11015\ : SRMux
    port map (
            O => \N__47011\,
            I => \N__46662\
        );

    \I__11014\ : SRMux
    port map (
            O => \N__47010\,
            I => \N__46662\
        );

    \I__11013\ : SRMux
    port map (
            O => \N__47009\,
            I => \N__46662\
        );

    \I__11012\ : SRMux
    port map (
            O => \N__47008\,
            I => \N__46662\
        );

    \I__11011\ : SRMux
    port map (
            O => \N__47007\,
            I => \N__46662\
        );

    \I__11010\ : SRMux
    port map (
            O => \N__47006\,
            I => \N__46662\
        );

    \I__11009\ : SRMux
    port map (
            O => \N__47005\,
            I => \N__46662\
        );

    \I__11008\ : SRMux
    port map (
            O => \N__47004\,
            I => \N__46662\
        );

    \I__11007\ : SRMux
    port map (
            O => \N__47003\,
            I => \N__46662\
        );

    \I__11006\ : SRMux
    port map (
            O => \N__47002\,
            I => \N__46662\
        );

    \I__11005\ : SRMux
    port map (
            O => \N__47001\,
            I => \N__46662\
        );

    \I__11004\ : SRMux
    port map (
            O => \N__47000\,
            I => \N__46662\
        );

    \I__11003\ : SRMux
    port map (
            O => \N__46999\,
            I => \N__46662\
        );

    \I__11002\ : SRMux
    port map (
            O => \N__46998\,
            I => \N__46662\
        );

    \I__11001\ : SRMux
    port map (
            O => \N__46997\,
            I => \N__46662\
        );

    \I__11000\ : SRMux
    port map (
            O => \N__46996\,
            I => \N__46662\
        );

    \I__10999\ : SRMux
    port map (
            O => \N__46995\,
            I => \N__46662\
        );

    \I__10998\ : SRMux
    port map (
            O => \N__46994\,
            I => \N__46662\
        );

    \I__10997\ : SRMux
    port map (
            O => \N__46993\,
            I => \N__46662\
        );

    \I__10996\ : SRMux
    port map (
            O => \N__46992\,
            I => \N__46662\
        );

    \I__10995\ : SRMux
    port map (
            O => \N__46991\,
            I => \N__46662\
        );

    \I__10994\ : SRMux
    port map (
            O => \N__46990\,
            I => \N__46662\
        );

    \I__10993\ : SRMux
    port map (
            O => \N__46989\,
            I => \N__46662\
        );

    \I__10992\ : SRMux
    port map (
            O => \N__46988\,
            I => \N__46662\
        );

    \I__10991\ : SRMux
    port map (
            O => \N__46987\,
            I => \N__46662\
        );

    \I__10990\ : SRMux
    port map (
            O => \N__46986\,
            I => \N__46662\
        );

    \I__10989\ : SRMux
    port map (
            O => \N__46985\,
            I => \N__46662\
        );

    \I__10988\ : SRMux
    port map (
            O => \N__46984\,
            I => \N__46662\
        );

    \I__10987\ : SRMux
    port map (
            O => \N__46983\,
            I => \N__46662\
        );

    \I__10986\ : SRMux
    port map (
            O => \N__46982\,
            I => \N__46662\
        );

    \I__10985\ : SRMux
    port map (
            O => \N__46981\,
            I => \N__46662\
        );

    \I__10984\ : SRMux
    port map (
            O => \N__46980\,
            I => \N__46662\
        );

    \I__10983\ : SRMux
    port map (
            O => \N__46979\,
            I => \N__46662\
        );

    \I__10982\ : SRMux
    port map (
            O => \N__46978\,
            I => \N__46662\
        );

    \I__10981\ : SRMux
    port map (
            O => \N__46977\,
            I => \N__46662\
        );

    \I__10980\ : SRMux
    port map (
            O => \N__46976\,
            I => \N__46662\
        );

    \I__10979\ : SRMux
    port map (
            O => \N__46975\,
            I => \N__46662\
        );

    \I__10978\ : SRMux
    port map (
            O => \N__46974\,
            I => \N__46662\
        );

    \I__10977\ : SRMux
    port map (
            O => \N__46973\,
            I => \N__46662\
        );

    \I__10976\ : SRMux
    port map (
            O => \N__46972\,
            I => \N__46662\
        );

    \I__10975\ : SRMux
    port map (
            O => \N__46971\,
            I => \N__46662\
        );

    \I__10974\ : SRMux
    port map (
            O => \N__46970\,
            I => \N__46662\
        );

    \I__10973\ : SRMux
    port map (
            O => \N__46969\,
            I => \N__46662\
        );

    \I__10972\ : SRMux
    port map (
            O => \N__46968\,
            I => \N__46662\
        );

    \I__10971\ : SRMux
    port map (
            O => \N__46967\,
            I => \N__46662\
        );

    \I__10970\ : SRMux
    port map (
            O => \N__46966\,
            I => \N__46662\
        );

    \I__10969\ : SRMux
    port map (
            O => \N__46965\,
            I => \N__46662\
        );

    \I__10968\ : SRMux
    port map (
            O => \N__46964\,
            I => \N__46662\
        );

    \I__10967\ : SRMux
    port map (
            O => \N__46963\,
            I => \N__46662\
        );

    \I__10966\ : SRMux
    port map (
            O => \N__46962\,
            I => \N__46662\
        );

    \I__10965\ : SRMux
    port map (
            O => \N__46961\,
            I => \N__46662\
        );

    \I__10964\ : SRMux
    port map (
            O => \N__46960\,
            I => \N__46662\
        );

    \I__10963\ : SRMux
    port map (
            O => \N__46959\,
            I => \N__46662\
        );

    \I__10962\ : SRMux
    port map (
            O => \N__46958\,
            I => \N__46662\
        );

    \I__10961\ : SRMux
    port map (
            O => \N__46957\,
            I => \N__46662\
        );

    \I__10960\ : SRMux
    port map (
            O => \N__46956\,
            I => \N__46662\
        );

    \I__10959\ : SRMux
    port map (
            O => \N__46955\,
            I => \N__46662\
        );

    \I__10958\ : GlobalMux
    port map (
            O => \N__46662\,
            I => \N__46659\
        );

    \I__10957\ : gio2CtrlBuf
    port map (
            O => \N__46659\,
            I => red_c_g
        );

    \I__10956\ : CascadeMux
    port map (
            O => \N__46656\,
            I => \N__46652\
        );

    \I__10955\ : InMux
    port map (
            O => \N__46655\,
            I => \N__46647\
        );

    \I__10954\ : InMux
    port map (
            O => \N__46652\,
            I => \N__46644\
        );

    \I__10953\ : InMux
    port map (
            O => \N__46651\,
            I => \N__46641\
        );

    \I__10952\ : InMux
    port map (
            O => \N__46650\,
            I => \N__46638\
        );

    \I__10951\ : LocalMux
    port map (
            O => \N__46647\,
            I => \N__46634\
        );

    \I__10950\ : LocalMux
    port map (
            O => \N__46644\,
            I => \N__46631\
        );

    \I__10949\ : LocalMux
    port map (
            O => \N__46641\,
            I => \N__46626\
        );

    \I__10948\ : LocalMux
    port map (
            O => \N__46638\,
            I => \N__46626\
        );

    \I__10947\ : InMux
    port map (
            O => \N__46637\,
            I => \N__46623\
        );

    \I__10946\ : Span4Mux_h
    port map (
            O => \N__46634\,
            I => \N__46620\
        );

    \I__10945\ : Span4Mux_h
    port map (
            O => \N__46631\,
            I => \N__46613\
        );

    \I__10944\ : Span4Mux_v
    port map (
            O => \N__46626\,
            I => \N__46613\
        );

    \I__10943\ : LocalMux
    port map (
            O => \N__46623\,
            I => \N__46613\
        );

    \I__10942\ : Odrv4
    port map (
            O => \N__46620\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10941\ : Odrv4
    port map (
            O => \N__46613\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__10940\ : CascadeMux
    port map (
            O => \N__46608\,
            I => \N__46605\
        );

    \I__10939\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46601\
        );

    \I__10938\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46598\
        );

    \I__10937\ : LocalMux
    port map (
            O => \N__46601\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__10936\ : LocalMux
    port map (
            O => \N__46598\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__10935\ : InMux
    port map (
            O => \N__46593\,
            I => \N__46589\
        );

    \I__10934\ : CascadeMux
    port map (
            O => \N__46592\,
            I => \N__46584\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__46589\,
            I => \N__46581\
        );

    \I__10932\ : InMux
    port map (
            O => \N__46588\,
            I => \N__46578\
        );

    \I__10931\ : InMux
    port map (
            O => \N__46587\,
            I => \N__46573\
        );

    \I__10930\ : InMux
    port map (
            O => \N__46584\,
            I => \N__46573\
        );

    \I__10929\ : Span4Mux_v
    port map (
            O => \N__46581\,
            I => \N__46568\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__46578\,
            I => \N__46568\
        );

    \I__10927\ : LocalMux
    port map (
            O => \N__46573\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10926\ : Odrv4
    port map (
            O => \N__46568\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__10925\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46560\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__46560\,
            I => \N__46555\
        );

    \I__10923\ : InMux
    port map (
            O => \N__46559\,
            I => \N__46550\
        );

    \I__10922\ : InMux
    port map (
            O => \N__46558\,
            I => \N__46550\
        );

    \I__10921\ : Span4Mux_v
    port map (
            O => \N__46555\,
            I => \N__46547\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__46550\,
            I => \N__46543\
        );

    \I__10919\ : Sp12to4
    port map (
            O => \N__46547\,
            I => \N__46540\
        );

    \I__10918\ : InMux
    port map (
            O => \N__46546\,
            I => \N__46537\
        );

    \I__10917\ : Span4Mux_v
    port map (
            O => \N__46543\,
            I => \N__46533\
        );

    \I__10916\ : Span12Mux_h
    port map (
            O => \N__46540\,
            I => \N__46530\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__46537\,
            I => \N__46527\
        );

    \I__10914\ : InMux
    port map (
            O => \N__46536\,
            I => \N__46524\
        );

    \I__10913\ : Span4Mux_h
    port map (
            O => \N__46533\,
            I => \N__46521\
        );

    \I__10912\ : Odrv12
    port map (
            O => \N__46530\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__10911\ : Odrv12
    port map (
            O => \N__46527\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__46524\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__10909\ : Odrv4
    port map (
            O => \N__46521\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__10908\ : CascadeMux
    port map (
            O => \N__46512\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\
        );

    \I__10907\ : InMux
    port map (
            O => \N__46509\,
            I => \N__46506\
        );

    \I__10906\ : LocalMux
    port map (
            O => \N__46506\,
            I => \N__46503\
        );

    \I__10905\ : Span4Mux_v
    port map (
            O => \N__46503\,
            I => \N__46498\
        );

    \I__10904\ : InMux
    port map (
            O => \N__46502\,
            I => \N__46493\
        );

    \I__10903\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46493\
        );

    \I__10902\ : Sp12to4
    port map (
            O => \N__46498\,
            I => \N__46488\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__46493\,
            I => \N__46488\
        );

    \I__10900\ : Span12Mux_h
    port map (
            O => \N__46488\,
            I => \N__46484\
        );

    \I__10899\ : InMux
    port map (
            O => \N__46487\,
            I => \N__46481\
        );

    \I__10898\ : Odrv12
    port map (
            O => \N__46484\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10897\ : LocalMux
    port map (
            O => \N__46481\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__10896\ : InMux
    port map (
            O => \N__46476\,
            I => \N__46470\
        );

    \I__10895\ : InMux
    port map (
            O => \N__46475\,
            I => \N__46470\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__46470\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__10893\ : InMux
    port map (
            O => \N__46467\,
            I => \N__46463\
        );

    \I__10892\ : InMux
    port map (
            O => \N__46466\,
            I => \N__46460\
        );

    \I__10891\ : LocalMux
    port map (
            O => \N__46463\,
            I => \N__46457\
        );

    \I__10890\ : LocalMux
    port map (
            O => \N__46460\,
            I => \N__46452\
        );

    \I__10889\ : Span4Mux_h
    port map (
            O => \N__46457\,
            I => \N__46449\
        );

    \I__10888\ : InMux
    port map (
            O => \N__46456\,
            I => \N__46446\
        );

    \I__10887\ : InMux
    port map (
            O => \N__46455\,
            I => \N__46443\
        );

    \I__10886\ : Span4Mux_v
    port map (
            O => \N__46452\,
            I => \N__46440\
        );

    \I__10885\ : Sp12to4
    port map (
            O => \N__46449\,
            I => \N__46435\
        );

    \I__10884\ : LocalMux
    port map (
            O => \N__46446\,
            I => \N__46435\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__46443\,
            I => \N__46430\
        );

    \I__10882\ : Sp12to4
    port map (
            O => \N__46440\,
            I => \N__46425\
        );

    \I__10881\ : Span12Mux_s8_v
    port map (
            O => \N__46435\,
            I => \N__46425\
        );

    \I__10880\ : InMux
    port map (
            O => \N__46434\,
            I => \N__46420\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46433\,
            I => \N__46420\
        );

    \I__10878\ : Odrv12
    port map (
            O => \N__46430\,
            I => phase_controller_inst1_state_4
        );

    \I__10877\ : Odrv12
    port map (
            O => \N__46425\,
            I => phase_controller_inst1_state_4
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__46420\,
            I => phase_controller_inst1_state_4
        );

    \I__10875\ : InMux
    port map (
            O => \N__46413\,
            I => \N__46410\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46410\,
            I => \N__46407\
        );

    \I__10873\ : Span4Mux_v
    port map (
            O => \N__46407\,
            I => \N__46404\
        );

    \I__10872\ : Span4Mux_h
    port map (
            O => \N__46404\,
            I => \N__46401\
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__46401\,
            I => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\
        );

    \I__10870\ : InMux
    port map (
            O => \N__46398\,
            I => \N__46395\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__46395\,
            I => \N__46392\
        );

    \I__10868\ : Span4Mux_h
    port map (
            O => \N__46392\,
            I => \N__46389\
        );

    \I__10867\ : Span4Mux_h
    port map (
            O => \N__46389\,
            I => \N__46385\
        );

    \I__10866\ : InMux
    port map (
            O => \N__46388\,
            I => \N__46382\
        );

    \I__10865\ : Odrv4
    port map (
            O => \N__46385\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__10864\ : LocalMux
    port map (
            O => \N__46382\,
            I => \phase_controller_inst1.state_RNI7NN7Z0Z_0\
        );

    \I__10863\ : CascadeMux
    port map (
            O => \N__46377\,
            I => \N__46374\
        );

    \I__10862\ : InMux
    port map (
            O => \N__46374\,
            I => \N__46369\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46366\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46372\,
            I => \N__46363\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__46369\,
            I => \N__46360\
        );

    \I__10858\ : LocalMux
    port map (
            O => \N__46366\,
            I => \N__46357\
        );

    \I__10857\ : LocalMux
    port map (
            O => \N__46363\,
            I => \N__46354\
        );

    \I__10856\ : Span4Mux_h
    port map (
            O => \N__46360\,
            I => \N__46350\
        );

    \I__10855\ : Span4Mux_h
    port map (
            O => \N__46357\,
            I => \N__46345\
        );

    \I__10854\ : Span4Mux_v
    port map (
            O => \N__46354\,
            I => \N__46345\
        );

    \I__10853\ : InMux
    port map (
            O => \N__46353\,
            I => \N__46342\
        );

    \I__10852\ : Odrv4
    port map (
            O => \N__46350\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10851\ : Odrv4
    port map (
            O => \N__46345\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10850\ : LocalMux
    port map (
            O => \N__46342\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__10849\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46332\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46329\
        );

    \I__10847\ : Span4Mux_h
    port map (
            O => \N__46329\,
            I => \N__46326\
        );

    \I__10846\ : Odrv4
    port map (
            O => \N__46326\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__10845\ : CascadeMux
    port map (
            O => \N__46323\,
            I => \N__46320\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46320\,
            I => \N__46315\
        );

    \I__10843\ : InMux
    port map (
            O => \N__46319\,
            I => \N__46312\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46318\,
            I => \N__46309\
        );

    \I__10841\ : LocalMux
    port map (
            O => \N__46315\,
            I => \N__46304\
        );

    \I__10840\ : LocalMux
    port map (
            O => \N__46312\,
            I => \N__46304\
        );

    \I__10839\ : LocalMux
    port map (
            O => \N__46309\,
            I => \N__46301\
        );

    \I__10838\ : Span4Mux_v
    port map (
            O => \N__46304\,
            I => \N__46295\
        );

    \I__10837\ : Span4Mux_v
    port map (
            O => \N__46301\,
            I => \N__46295\
        );

    \I__10836\ : InMux
    port map (
            O => \N__46300\,
            I => \N__46292\
        );

    \I__10835\ : Odrv4
    port map (
            O => \N__46295\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__46292\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46287\,
            I => \N__46284\
        );

    \I__10832\ : LocalMux
    port map (
            O => \N__46284\,
            I => \N__46281\
        );

    \I__10831\ : Span4Mux_h
    port map (
            O => \N__46281\,
            I => \N__46278\
        );

    \I__10830\ : Odrv4
    port map (
            O => \N__46278\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__10829\ : CascadeMux
    port map (
            O => \N__46275\,
            I => \N__46272\
        );

    \I__10828\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46268\
        );

    \I__10827\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46264\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__46268\,
            I => \N__46261\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46267\,
            I => \N__46258\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__46264\,
            I => \N__46255\
        );

    \I__10823\ : Span4Mux_v
    port map (
            O => \N__46261\,
            I => \N__46252\
        );

    \I__10822\ : LocalMux
    port map (
            O => \N__46258\,
            I => \N__46249\
        );

    \I__10821\ : Span4Mux_h
    port map (
            O => \N__46255\,
            I => \N__46245\
        );

    \I__10820\ : Span4Mux_h
    port map (
            O => \N__46252\,
            I => \N__46240\
        );

    \I__10819\ : Span4Mux_v
    port map (
            O => \N__46249\,
            I => \N__46240\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46248\,
            I => \N__46237\
        );

    \I__10817\ : Odrv4
    port map (
            O => \N__46245\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10816\ : Odrv4
    port map (
            O => \N__46240\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46237\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46230\,
            I => \N__46227\
        );

    \I__10813\ : LocalMux
    port map (
            O => \N__46227\,
            I => \N__46224\
        );

    \I__10812\ : Span4Mux_h
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__10811\ : Odrv4
    port map (
            O => \N__46221\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__10810\ : InMux
    port map (
            O => \N__46218\,
            I => \N__46214\
        );

    \I__10809\ : InMux
    port map (
            O => \N__46217\,
            I => \N__46211\
        );

    \I__10808\ : LocalMux
    port map (
            O => \N__46214\,
            I => \N__46205\
        );

    \I__10807\ : LocalMux
    port map (
            O => \N__46211\,
            I => \N__46205\
        );

    \I__10806\ : InMux
    port map (
            O => \N__46210\,
            I => \N__46201\
        );

    \I__10805\ : Span4Mux_v
    port map (
            O => \N__46205\,
            I => \N__46198\
        );

    \I__10804\ : InMux
    port map (
            O => \N__46204\,
            I => \N__46195\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__46201\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10802\ : Odrv4
    port map (
            O => \N__46198\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46195\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__10800\ : InMux
    port map (
            O => \N__46188\,
            I => \N__46185\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__46185\,
            I => \N__46182\
        );

    \I__10798\ : Span4Mux_h
    port map (
            O => \N__46182\,
            I => \N__46179\
        );

    \I__10797\ : Odrv4
    port map (
            O => \N__46179\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__10796\ : InMux
    port map (
            O => \N__46176\,
            I => \N__46173\
        );

    \I__10795\ : LocalMux
    port map (
            O => \N__46173\,
            I => \N__46168\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46172\,
            I => \N__46165\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46171\,
            I => \N__46162\
        );

    \I__10792\ : Span12Mux_s11_v
    port map (
            O => \N__46168\,
            I => \N__46157\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__46165\,
            I => \N__46157\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46162\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__10789\ : Odrv12
    port map (
            O => \N__46157\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46152\,
            I => \N__46149\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46143\
        );

    \I__10786\ : InMux
    port map (
            O => \N__46148\,
            I => \N__46140\
        );

    \I__10785\ : CascadeMux
    port map (
            O => \N__46147\,
            I => \N__46137\
        );

    \I__10784\ : InMux
    port map (
            O => \N__46146\,
            I => \N__46134\
        );

    \I__10783\ : Span4Mux_h
    port map (
            O => \N__46143\,
            I => \N__46131\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__46140\,
            I => \N__46128\
        );

    \I__10781\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46125\
        );

    \I__10780\ : LocalMux
    port map (
            O => \N__46134\,
            I => \N__46122\
        );

    \I__10779\ : Span4Mux_h
    port map (
            O => \N__46131\,
            I => \N__46117\
        );

    \I__10778\ : Span4Mux_v
    port map (
            O => \N__46128\,
            I => \N__46117\
        );

    \I__10777\ : LocalMux
    port map (
            O => \N__46125\,
            I => \N__46114\
        );

    \I__10776\ : Odrv12
    port map (
            O => \N__46122\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__46117\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__10774\ : Odrv4
    port map (
            O => \N__46114\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__10773\ : InMux
    port map (
            O => \N__46107\,
            I => \N__46104\
        );

    \I__10772\ : LocalMux
    port map (
            O => \N__46104\,
            I => \N__46101\
        );

    \I__10771\ : Span4Mux_h
    port map (
            O => \N__46101\,
            I => \N__46098\
        );

    \I__10770\ : Odrv4
    port map (
            O => \N__46098\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46095\,
            I => \N__46092\
        );

    \I__10768\ : LocalMux
    port map (
            O => \N__46092\,
            I => \N__46089\
        );

    \I__10767\ : Span4Mux_h
    port map (
            O => \N__46089\,
            I => \N__46086\
        );

    \I__10766\ : Odrv4
    port map (
            O => \N__46086\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__10765\ : CEMux
    port map (
            O => \N__46083\,
            I => \N__46059\
        );

    \I__10764\ : CEMux
    port map (
            O => \N__46082\,
            I => \N__46059\
        );

    \I__10763\ : CEMux
    port map (
            O => \N__46081\,
            I => \N__46059\
        );

    \I__10762\ : CEMux
    port map (
            O => \N__46080\,
            I => \N__46059\
        );

    \I__10761\ : CEMux
    port map (
            O => \N__46079\,
            I => \N__46059\
        );

    \I__10760\ : CEMux
    port map (
            O => \N__46078\,
            I => \N__46059\
        );

    \I__10759\ : CEMux
    port map (
            O => \N__46077\,
            I => \N__46059\
        );

    \I__10758\ : CEMux
    port map (
            O => \N__46076\,
            I => \N__46059\
        );

    \I__10757\ : GlobalMux
    port map (
            O => \N__46059\,
            I => \N__46056\
        );

    \I__10756\ : gio2CtrlBuf
    port map (
            O => \N__46056\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__10755\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46050\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__46050\,
            I => \N__46047\
        );

    \I__10753\ : Odrv12
    port map (
            O => \N__46047\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46044\,
            I => \N__46038\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46043\,
            I => \N__46038\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46038\,
            I => \N__46034\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46031\
        );

    \I__10748\ : Span4Mux_h
    port map (
            O => \N__46034\,
            I => \N__46028\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__46031\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10746\ : Odrv4
    port map (
            O => \N__46028\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10745\ : CascadeMux
    port map (
            O => \N__46023\,
            I => \N__46019\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46022\,
            I => \N__46014\
        );

    \I__10743\ : InMux
    port map (
            O => \N__46019\,
            I => \N__46014\
        );

    \I__10742\ : LocalMux
    port map (
            O => \N__46014\,
            I => \N__46010\
        );

    \I__10741\ : InMux
    port map (
            O => \N__46013\,
            I => \N__46007\
        );

    \I__10740\ : Span4Mux_h
    port map (
            O => \N__46010\,
            I => \N__46004\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46007\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__46004\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10737\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45993\
        );

    \I__10736\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45993\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__45993\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__10734\ : CascadeMux
    port map (
            O => \N__45990\,
            I => \N__45987\
        );

    \I__10733\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45984\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__45984\,
            I => \N__45981\
        );

    \I__10731\ : Odrv12
    port map (
            O => \N__45981\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__10730\ : CascadeMux
    port map (
            O => \N__45978\,
            I => \N__45974\
        );

    \I__10729\ : InMux
    port map (
            O => \N__45977\,
            I => \N__45971\
        );

    \I__10728\ : InMux
    port map (
            O => \N__45974\,
            I => \N__45968\
        );

    \I__10727\ : LocalMux
    port map (
            O => \N__45971\,
            I => \N__45963\
        );

    \I__10726\ : LocalMux
    port map (
            O => \N__45968\,
            I => \N__45963\
        );

    \I__10725\ : Span4Mux_v
    port map (
            O => \N__45963\,
            I => \N__45960\
        );

    \I__10724\ : Odrv4
    port map (
            O => \N__45960\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__10723\ : InMux
    port map (
            O => \N__45957\,
            I => \N__45954\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__45954\,
            I => \N__45950\
        );

    \I__10721\ : InMux
    port map (
            O => \N__45953\,
            I => \N__45946\
        );

    \I__10720\ : Span4Mux_h
    port map (
            O => \N__45950\,
            I => \N__45943\
        );

    \I__10719\ : InMux
    port map (
            O => \N__45949\,
            I => \N__45940\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__45946\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10717\ : Odrv4
    port map (
            O => \N__45943\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__45940\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10715\ : CascadeMux
    port map (
            O => \N__45933\,
            I => \N__45930\
        );

    \I__10714\ : InMux
    port map (
            O => \N__45930\,
            I => \N__45927\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__45927\,
            I => \N__45922\
        );

    \I__10712\ : InMux
    port map (
            O => \N__45926\,
            I => \N__45919\
        );

    \I__10711\ : InMux
    port map (
            O => \N__45925\,
            I => \N__45916\
        );

    \I__10710\ : Span4Mux_v
    port map (
            O => \N__45922\,
            I => \N__45913\
        );

    \I__10709\ : LocalMux
    port map (
            O => \N__45919\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__45916\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__45913\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10706\ : InMux
    port map (
            O => \N__45906\,
            I => \N__45902\
        );

    \I__10705\ : InMux
    port map (
            O => \N__45905\,
            I => \N__45899\
        );

    \I__10704\ : LocalMux
    port map (
            O => \N__45902\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__10703\ : LocalMux
    port map (
            O => \N__45899\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__10702\ : CascadeMux
    port map (
            O => \N__45894\,
            I => \N__45891\
        );

    \I__10701\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45888\
        );

    \I__10700\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45885\
        );

    \I__10699\ : Odrv12
    port map (
            O => \N__45885\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__10698\ : CascadeMux
    port map (
            O => \N__45882\,
            I => \N__45879\
        );

    \I__10697\ : InMux
    port map (
            O => \N__45879\,
            I => \N__45876\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__45876\,
            I => \N__45873\
        );

    \I__10695\ : Span4Mux_v
    port map (
            O => \N__45873\,
            I => \N__45870\
        );

    \I__10694\ : Span4Mux_h
    port map (
            O => \N__45870\,
            I => \N__45867\
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__45867\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__10692\ : CascadeMux
    port map (
            O => \N__45864\,
            I => \N__45860\
        );

    \I__10691\ : InMux
    port map (
            O => \N__45863\,
            I => \N__45855\
        );

    \I__10690\ : InMux
    port map (
            O => \N__45860\,
            I => \N__45855\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__45855\,
            I => \N__45851\
        );

    \I__10688\ : InMux
    port map (
            O => \N__45854\,
            I => \N__45848\
        );

    \I__10687\ : Span4Mux_h
    port map (
            O => \N__45851\,
            I => \N__45845\
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__45848\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10685\ : Odrv4
    port map (
            O => \N__45845\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10684\ : CascadeMux
    port map (
            O => \N__45840\,
            I => \N__45836\
        );

    \I__10683\ : InMux
    port map (
            O => \N__45839\,
            I => \N__45832\
        );

    \I__10682\ : InMux
    port map (
            O => \N__45836\,
            I => \N__45827\
        );

    \I__10681\ : InMux
    port map (
            O => \N__45835\,
            I => \N__45827\
        );

    \I__10680\ : LocalMux
    port map (
            O => \N__45832\,
            I => \N__45822\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__45827\,
            I => \N__45822\
        );

    \I__10678\ : Odrv4
    port map (
            O => \N__45822\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10677\ : InMux
    port map (
            O => \N__45819\,
            I => \N__45816\
        );

    \I__10676\ : LocalMux
    port map (
            O => \N__45816\,
            I => \N__45813\
        );

    \I__10675\ : Span4Mux_v
    port map (
            O => \N__45813\,
            I => \N__45810\
        );

    \I__10674\ : Span4Mux_h
    port map (
            O => \N__45810\,
            I => \N__45807\
        );

    \I__10673\ : Odrv4
    port map (
            O => \N__45807\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__10672\ : InMux
    port map (
            O => \N__45804\,
            I => \N__45801\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__45801\,
            I => \N__45797\
        );

    \I__10670\ : InMux
    port map (
            O => \N__45800\,
            I => \N__45794\
        );

    \I__10669\ : Odrv4
    port map (
            O => \N__45797\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__45794\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__10667\ : CascadeMux
    port map (
            O => \N__45789\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\
        );

    \I__10666\ : InMux
    port map (
            O => \N__45786\,
            I => \N__45783\
        );

    \I__10665\ : LocalMux
    port map (
            O => \N__45783\,
            I => \N__45778\
        );

    \I__10664\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45773\
        );

    \I__10663\ : InMux
    port map (
            O => \N__45781\,
            I => \N__45773\
        );

    \I__10662\ : Span4Mux_h
    port map (
            O => \N__45778\,
            I => \N__45768\
        );

    \I__10661\ : LocalMux
    port map (
            O => \N__45773\,
            I => \N__45768\
        );

    \I__10660\ : Span4Mux_v
    port map (
            O => \N__45768\,
            I => \N__45764\
        );

    \I__10659\ : CascadeMux
    port map (
            O => \N__45767\,
            I => \N__45761\
        );

    \I__10658\ : Span4Mux_h
    port map (
            O => \N__45764\,
            I => \N__45758\
        );

    \I__10657\ : InMux
    port map (
            O => \N__45761\,
            I => \N__45755\
        );

    \I__10656\ : Odrv4
    port map (
            O => \N__45758\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__45755\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__10654\ : InMux
    port map (
            O => \N__45750\,
            I => \N__45744\
        );

    \I__10653\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45744\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__45744\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__10651\ : InMux
    port map (
            O => \N__45741\,
            I => \N__45738\
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__45738\,
            I => \N__45734\
        );

    \I__10649\ : InMux
    port map (
            O => \N__45737\,
            I => \N__45731\
        );

    \I__10648\ : Odrv4
    port map (
            O => \N__45734\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10647\ : LocalMux
    port map (
            O => \N__45731\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__10646\ : InMux
    port map (
            O => \N__45726\,
            I => \N__45720\
        );

    \I__10645\ : InMux
    port map (
            O => \N__45725\,
            I => \N__45720\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__45720\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__10643\ : InMux
    port map (
            O => \N__45717\,
            I => \N__45711\
        );

    \I__10642\ : InMux
    port map (
            O => \N__45716\,
            I => \N__45711\
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__45711\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__10640\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45702\
        );

    \I__10639\ : InMux
    port map (
            O => \N__45707\,
            I => \N__45702\
        );

    \I__10638\ : LocalMux
    port map (
            O => \N__45702\,
            I => \N__45699\
        );

    \I__10637\ : Odrv4
    port map (
            O => \N__45699\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__10636\ : CascadeMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__10635\ : InMux
    port map (
            O => \N__45693\,
            I => \N__45687\
        );

    \I__10634\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45687\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__45687\,
            I => \N__45684\
        );

    \I__10632\ : Odrv4
    port map (
            O => \N__45684\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__10631\ : CascadeMux
    port map (
            O => \N__45681\,
            I => \N__45678\
        );

    \I__10630\ : InMux
    port map (
            O => \N__45678\,
            I => \N__45672\
        );

    \I__10629\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45672\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__45672\,
            I => \N__45669\
        );

    \I__10627\ : Odrv4
    port map (
            O => \N__45669\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__10626\ : InMux
    port map (
            O => \N__45666\,
            I => \N__45662\
        );

    \I__10625\ : InMux
    port map (
            O => \N__45665\,
            I => \N__45659\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__45662\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__45659\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__10622\ : CascadeMux
    port map (
            O => \N__45654\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__10621\ : InMux
    port map (
            O => \N__45651\,
            I => \N__45645\
        );

    \I__10620\ : InMux
    port map (
            O => \N__45650\,
            I => \N__45640\
        );

    \I__10619\ : InMux
    port map (
            O => \N__45649\,
            I => \N__45640\
        );

    \I__10618\ : InMux
    port map (
            O => \N__45648\,
            I => \N__45637\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__45645\,
            I => \N__45632\
        );

    \I__10616\ : LocalMux
    port map (
            O => \N__45640\,
            I => \N__45632\
        );

    \I__10615\ : LocalMux
    port map (
            O => \N__45637\,
            I => \N__45629\
        );

    \I__10614\ : Span4Mux_v
    port map (
            O => \N__45632\,
            I => \N__45626\
        );

    \I__10613\ : Span4Mux_h
    port map (
            O => \N__45629\,
            I => \N__45623\
        );

    \I__10612\ : Span4Mux_h
    port map (
            O => \N__45626\,
            I => \N__45620\
        );

    \I__10611\ : Span4Mux_h
    port map (
            O => \N__45623\,
            I => \N__45617\
        );

    \I__10610\ : Odrv4
    port map (
            O => \N__45620\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10609\ : Odrv4
    port map (
            O => \N__45617\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__10608\ : InMux
    port map (
            O => \N__45612\,
            I => \N__45608\
        );

    \I__10607\ : InMux
    port map (
            O => \N__45611\,
            I => \N__45605\
        );

    \I__10606\ : LocalMux
    port map (
            O => \N__45608\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__45605\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__10604\ : CascadeMux
    port map (
            O => \N__45600\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\
        );

    \I__10603\ : InMux
    port map (
            O => \N__45597\,
            I => \N__45592\
        );

    \I__10602\ : InMux
    port map (
            O => \N__45596\,
            I => \N__45587\
        );

    \I__10601\ : InMux
    port map (
            O => \N__45595\,
            I => \N__45587\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__45592\,
            I => \N__45581\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__45587\,
            I => \N__45581\
        );

    \I__10598\ : InMux
    port map (
            O => \N__45586\,
            I => \N__45578\
        );

    \I__10597\ : Span4Mux_v
    port map (
            O => \N__45581\,
            I => \N__45575\
        );

    \I__10596\ : LocalMux
    port map (
            O => \N__45578\,
            I => \N__45572\
        );

    \I__10595\ : Span4Mux_h
    port map (
            O => \N__45575\,
            I => \N__45569\
        );

    \I__10594\ : Span12Mux_h
    port map (
            O => \N__45572\,
            I => \N__45566\
        );

    \I__10593\ : Odrv4
    port map (
            O => \N__45569\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10592\ : Odrv12
    port map (
            O => \N__45566\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__10591\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45558\
        );

    \I__10590\ : LocalMux
    port map (
            O => \N__45558\,
            I => \N__45554\
        );

    \I__10589\ : InMux
    port map (
            O => \N__45557\,
            I => \N__45551\
        );

    \I__10588\ : Odrv4
    port map (
            O => \N__45554\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__45551\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__10586\ : CascadeMux
    port map (
            O => \N__45546\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\
        );

    \I__10585\ : InMux
    port map (
            O => \N__45543\,
            I => \N__45538\
        );

    \I__10584\ : InMux
    port map (
            O => \N__45542\,
            I => \N__45533\
        );

    \I__10583\ : InMux
    port map (
            O => \N__45541\,
            I => \N__45533\
        );

    \I__10582\ : LocalMux
    port map (
            O => \N__45538\,
            I => \N__45530\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__45533\,
            I => \N__45527\
        );

    \I__10580\ : Span4Mux_h
    port map (
            O => \N__45530\,
            I => \N__45524\
        );

    \I__10579\ : Span4Mux_h
    port map (
            O => \N__45527\,
            I => \N__45521\
        );

    \I__10578\ : Span4Mux_h
    port map (
            O => \N__45524\,
            I => \N__45517\
        );

    \I__10577\ : Span4Mux_h
    port map (
            O => \N__45521\,
            I => \N__45514\
        );

    \I__10576\ : InMux
    port map (
            O => \N__45520\,
            I => \N__45511\
        );

    \I__10575\ : Odrv4
    port map (
            O => \N__45517\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10574\ : Odrv4
    port map (
            O => \N__45514\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10573\ : LocalMux
    port map (
            O => \N__45511\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__10572\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45501\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__45501\,
            I => \N__45498\
        );

    \I__10570\ : Odrv4
    port map (
            O => \N__45498\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__10569\ : InMux
    port map (
            O => \N__45495\,
            I => \N__45490\
        );

    \I__10568\ : InMux
    port map (
            O => \N__45494\,
            I => \N__45485\
        );

    \I__10567\ : InMux
    port map (
            O => \N__45493\,
            I => \N__45485\
        );

    \I__10566\ : LocalMux
    port map (
            O => \N__45490\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__45485\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__10564\ : CascadeMux
    port map (
            O => \N__45480\,
            I => \N__45475\
        );

    \I__10563\ : InMux
    port map (
            O => \N__45479\,
            I => \N__45472\
        );

    \I__10562\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45467\
        );

    \I__10561\ : InMux
    port map (
            O => \N__45475\,
            I => \N__45467\
        );

    \I__10560\ : LocalMux
    port map (
            O => \N__45472\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10559\ : LocalMux
    port map (
            O => \N__45467\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45462\,
            I => \N__45456\
        );

    \I__10557\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45456\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__45456\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__10555\ : CascadeMux
    port map (
            O => \N__45453\,
            I => \N__45450\
        );

    \I__10554\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45447\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__45447\,
            I => \N__45444\
        );

    \I__10552\ : Odrv4
    port map (
            O => \N__45444\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__10551\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45438\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__45438\,
            I => \N__45435\
        );

    \I__10549\ : Span4Mux_v
    port map (
            O => \N__45435\,
            I => \N__45432\
        );

    \I__10548\ : Odrv4
    port map (
            O => \N__45432\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__45429\,
            I => \N__45424\
        );

    \I__10546\ : InMux
    port map (
            O => \N__45428\,
            I => \N__45421\
        );

    \I__10545\ : InMux
    port map (
            O => \N__45427\,
            I => \N__45416\
        );

    \I__10544\ : InMux
    port map (
            O => \N__45424\,
            I => \N__45416\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__45421\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45416\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__10541\ : CascadeMux
    port map (
            O => \N__45411\,
            I => \N__45406\
        );

    \I__10540\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45403\
        );

    \I__10539\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45398\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45398\
        );

    \I__10537\ : LocalMux
    port map (
            O => \N__45403\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__45398\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__10535\ : CascadeMux
    port map (
            O => \N__45393\,
            I => \N__45390\
        );

    \I__10534\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45387\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__45387\,
            I => \N__45384\
        );

    \I__10532\ : Span4Mux_v
    port map (
            O => \N__45384\,
            I => \N__45381\
        );

    \I__10531\ : Odrv4
    port map (
            O => \N__45381\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__10530\ : InMux
    port map (
            O => \N__45378\,
            I => \N__45374\
        );

    \I__10529\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45371\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__45374\,
            I => \N__45364\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__45371\,
            I => \N__45364\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45370\,
            I => \N__45361\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45369\,
            I => \N__45358\
        );

    \I__10524\ : Span12Mux_h
    port map (
            O => \N__45364\,
            I => \N__45355\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__45361\,
            I => \N__45350\
        );

    \I__10522\ : LocalMux
    port map (
            O => \N__45358\,
            I => \N__45350\
        );

    \I__10521\ : Odrv12
    port map (
            O => \N__45355\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10520\ : Odrv12
    port map (
            O => \N__45350\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45345\,
            I => \N__45341\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45344\,
            I => \N__45337\
        );

    \I__10517\ : LocalMux
    port map (
            O => \N__45341\,
            I => \N__45334\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45340\,
            I => \N__45331\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__45337\,
            I => \N__45326\
        );

    \I__10514\ : Span4Mux_h
    port map (
            O => \N__45334\,
            I => \N__45326\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__45331\,
            I => \N__45323\
        );

    \I__10512\ : Odrv4
    port map (
            O => \N__45326\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__10511\ : Odrv12
    port map (
            O => \N__45323\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45318\,
            I => \N__45313\
        );

    \I__10509\ : InMux
    port map (
            O => \N__45317\,
            I => \N__45310\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45316\,
            I => \N__45307\
        );

    \I__10507\ : LocalMux
    port map (
            O => \N__45313\,
            I => \N__45302\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__45310\,
            I => \N__45302\
        );

    \I__10505\ : LocalMux
    port map (
            O => \N__45307\,
            I => \N__45298\
        );

    \I__10504\ : Span4Mux_v
    port map (
            O => \N__45302\,
            I => \N__45295\
        );

    \I__10503\ : InMux
    port map (
            O => \N__45301\,
            I => \N__45292\
        );

    \I__10502\ : Span4Mux_h
    port map (
            O => \N__45298\,
            I => \N__45289\
        );

    \I__10501\ : Span4Mux_h
    port map (
            O => \N__45295\,
            I => \N__45284\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__45292\,
            I => \N__45284\
        );

    \I__10499\ : Odrv4
    port map (
            O => \N__45289\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10498\ : Odrv4
    port map (
            O => \N__45284\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__10497\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45276\
        );

    \I__10496\ : LocalMux
    port map (
            O => \N__45276\,
            I => \N__45272\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45275\,
            I => \N__45268\
        );

    \I__10494\ : Span4Mux_h
    port map (
            O => \N__45272\,
            I => \N__45265\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45271\,
            I => \N__45262\
        );

    \I__10492\ : LocalMux
    port map (
            O => \N__45268\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__10491\ : Odrv4
    port map (
            O => \N__45265\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45262\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__10489\ : InMux
    port map (
            O => \N__45255\,
            I => \N__45252\
        );

    \I__10488\ : LocalMux
    port map (
            O => \N__45252\,
            I => \N__45249\
        );

    \I__10487\ : Span4Mux_h
    port map (
            O => \N__45249\,
            I => \N__45246\
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__45246\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__10485\ : InMux
    port map (
            O => \N__45243\,
            I => \N__45238\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45233\
        );

    \I__10483\ : InMux
    port map (
            O => \N__45241\,
            I => \N__45233\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__45238\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__45233\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__10480\ : CascadeMux
    port map (
            O => \N__45228\,
            I => \N__45224\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45220\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45224\,
            I => \N__45215\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45223\,
            I => \N__45215\
        );

    \I__10476\ : LocalMux
    port map (
            O => \N__45220\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__45215\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__10474\ : CascadeMux
    port map (
            O => \N__45210\,
            I => \N__45207\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45207\,
            I => \N__45204\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45204\,
            I => \N__45201\
        );

    \I__10471\ : Span4Mux_h
    port map (
            O => \N__45201\,
            I => \N__45198\
        );

    \I__10470\ : Odrv4
    port map (
            O => \N__45198\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45195\,
            I => \N__45188\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45194\,
            I => \N__45188\
        );

    \I__10467\ : InMux
    port map (
            O => \N__45193\,
            I => \N__45185\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45188\,
            I => \N__45182\
        );

    \I__10465\ : LocalMux
    port map (
            O => \N__45185\,
            I => \N__45178\
        );

    \I__10464\ : Span4Mux_h
    port map (
            O => \N__45182\,
            I => \N__45175\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45181\,
            I => \N__45172\
        );

    \I__10462\ : Odrv12
    port map (
            O => \N__45178\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__45175\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__45172\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45165\,
            I => \N__45162\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45159\
        );

    \I__10457\ : Span4Mux_v
    port map (
            O => \N__45159\,
            I => \N__45155\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45158\,
            I => \N__45152\
        );

    \I__10455\ : Odrv4
    port map (
            O => \N__45155\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45152\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45141\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45141\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__45141\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45138\,
            I => \N__45135\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45135\,
            I => \N__45129\
        );

    \I__10448\ : InMux
    port map (
            O => \N__45134\,
            I => \N__45122\
        );

    \I__10447\ : InMux
    port map (
            O => \N__45133\,
            I => \N__45122\
        );

    \I__10446\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45122\
        );

    \I__10445\ : Odrv12
    port map (
            O => \N__45129\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10444\ : LocalMux
    port map (
            O => \N__45122\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45113\
        );

    \I__10442\ : CascadeMux
    port map (
            O => \N__45116\,
            I => \N__45110\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__45113\,
            I => \N__45107\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45110\,
            I => \N__45104\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__45107\,
            I => \N__45101\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__45104\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__45101\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__10436\ : CascadeMux
    port map (
            O => \N__45096\,
            I => \N__45093\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45093\,
            I => \N__45087\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45092\,
            I => \N__45087\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45087\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45084\,
            I => \N__45081\
        );

    \I__10431\ : LocalMux
    port map (
            O => \N__45081\,
            I => \N__45076\
        );

    \I__10430\ : InMux
    port map (
            O => \N__45080\,
            I => \N__45073\
        );

    \I__10429\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45070\
        );

    \I__10428\ : Span4Mux_h
    port map (
            O => \N__45076\,
            I => \N__45065\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45073\,
            I => \N__45065\
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45070\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__10425\ : Odrv4
    port map (
            O => \N__45065\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__10424\ : InMux
    port map (
            O => \N__45060\,
            I => \N__45057\
        );

    \I__10423\ : LocalMux
    port map (
            O => \N__45057\,
            I => \N__45053\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45056\,
            I => \N__45048\
        );

    \I__10421\ : Span4Mux_v
    port map (
            O => \N__45053\,
            I => \N__45045\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45052\,
            I => \N__45040\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45051\,
            I => \N__45040\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45048\,
            I => \N__45037\
        );

    \I__10417\ : Sp12to4
    port map (
            O => \N__45045\,
            I => \N__45032\
        );

    \I__10416\ : LocalMux
    port map (
            O => \N__45040\,
            I => \N__45032\
        );

    \I__10415\ : Odrv4
    port map (
            O => \N__45037\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__10414\ : Odrv12
    port map (
            O => \N__45032\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__10413\ : CascadeMux
    port map (
            O => \N__45027\,
            I => \N__45024\
        );

    \I__10412\ : InMux
    port map (
            O => \N__45024\,
            I => \N__45021\
        );

    \I__10411\ : LocalMux
    port map (
            O => \N__45021\,
            I => \N__45018\
        );

    \I__10410\ : Odrv4
    port map (
            O => \N__45018\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45015\,
            I => \N__45012\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__45012\,
            I => \N__45007\
        );

    \I__10407\ : InMux
    port map (
            O => \N__45011\,
            I => \N__45004\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45010\,
            I => \N__45001\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__45007\,
            I => \N__44996\
        );

    \I__10404\ : LocalMux
    port map (
            O => \N__45004\,
            I => \N__44996\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45001\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__10402\ : Odrv4
    port map (
            O => \N__44996\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__10401\ : InMux
    port map (
            O => \N__44991\,
            I => \N__44987\
        );

    \I__10400\ : InMux
    port map (
            O => \N__44990\,
            I => \N__44984\
        );

    \I__10399\ : LocalMux
    port map (
            O => \N__44987\,
            I => \N__44980\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__44984\,
            I => \N__44977\
        );

    \I__10397\ : InMux
    port map (
            O => \N__44983\,
            I => \N__44973\
        );

    \I__10396\ : Span4Mux_v
    port map (
            O => \N__44980\,
            I => \N__44968\
        );

    \I__10395\ : Span4Mux_v
    port map (
            O => \N__44977\,
            I => \N__44968\
        );

    \I__10394\ : InMux
    port map (
            O => \N__44976\,
            I => \N__44965\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__44973\,
            I => \N__44962\
        );

    \I__10392\ : Sp12to4
    port map (
            O => \N__44968\,
            I => \N__44957\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__44965\,
            I => \N__44957\
        );

    \I__10390\ : Odrv4
    port map (
            O => \N__44962\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__10389\ : Odrv12
    port map (
            O => \N__44957\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__10388\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44949\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44946\
        );

    \I__10386\ : Span4Mux_h
    port map (
            O => \N__44946\,
            I => \N__44943\
        );

    \I__10385\ : Odrv4
    port map (
            O => \N__44943\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__10384\ : InMux
    port map (
            O => \N__44940\,
            I => \N__44937\
        );

    \I__10383\ : LocalMux
    port map (
            O => \N__44937\,
            I => \N__44934\
        );

    \I__10382\ : Odrv4
    port map (
            O => \N__44934\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__10381\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44926\
        );

    \I__10380\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44921\
        );

    \I__10379\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44921\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__44926\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__44921\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__10376\ : CascadeMux
    port map (
            O => \N__44916\,
            I => \N__44911\
        );

    \I__10375\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44908\
        );

    \I__10374\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44903\
        );

    \I__10373\ : InMux
    port map (
            O => \N__44911\,
            I => \N__44903\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__44908\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10371\ : LocalMux
    port map (
            O => \N__44903\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__10370\ : CascadeMux
    port map (
            O => \N__44898\,
            I => \N__44895\
        );

    \I__10369\ : InMux
    port map (
            O => \N__44895\,
            I => \N__44892\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__44892\,
            I => \N__44889\
        );

    \I__10367\ : Odrv12
    port map (
            O => \N__44889\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__10366\ : InMux
    port map (
            O => \N__44886\,
            I => \N__44881\
        );

    \I__10365\ : InMux
    port map (
            O => \N__44885\,
            I => \N__44878\
        );

    \I__10364\ : InMux
    port map (
            O => \N__44884\,
            I => \N__44875\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__44881\,
            I => \N__44872\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__44878\,
            I => \N__44868\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__44875\,
            I => \N__44865\
        );

    \I__10360\ : Span4Mux_v
    port map (
            O => \N__44872\,
            I => \N__44862\
        );

    \I__10359\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44859\
        );

    \I__10358\ : Span4Mux_v
    port map (
            O => \N__44868\,
            I => \N__44852\
        );

    \I__10357\ : Span4Mux_v
    port map (
            O => \N__44865\,
            I => \N__44852\
        );

    \I__10356\ : Span4Mux_h
    port map (
            O => \N__44862\,
            I => \N__44852\
        );

    \I__10355\ : LocalMux
    port map (
            O => \N__44859\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__10354\ : Odrv4
    port map (
            O => \N__44852\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__10353\ : CascadeMux
    port map (
            O => \N__44847\,
            I => \N__44844\
        );

    \I__10352\ : InMux
    port map (
            O => \N__44844\,
            I => \N__44839\
        );

    \I__10351\ : InMux
    port map (
            O => \N__44843\,
            I => \N__44834\
        );

    \I__10350\ : InMux
    port map (
            O => \N__44842\,
            I => \N__44834\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__44839\,
            I => \N__44831\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__44834\,
            I => \N__44827\
        );

    \I__10347\ : Span4Mux_v
    port map (
            O => \N__44831\,
            I => \N__44824\
        );

    \I__10346\ : InMux
    port map (
            O => \N__44830\,
            I => \N__44821\
        );

    \I__10345\ : Span4Mux_h
    port map (
            O => \N__44827\,
            I => \N__44818\
        );

    \I__10344\ : Span4Mux_h
    port map (
            O => \N__44824\,
            I => \N__44815\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__44821\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__10342\ : Odrv4
    port map (
            O => \N__44818\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__10341\ : Odrv4
    port map (
            O => \N__44815\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__10340\ : InMux
    port map (
            O => \N__44808\,
            I => \N__44802\
        );

    \I__10339\ : InMux
    port map (
            O => \N__44807\,
            I => \N__44799\
        );

    \I__10338\ : InMux
    port map (
            O => \N__44806\,
            I => \N__44796\
        );

    \I__10337\ : InMux
    port map (
            O => \N__44805\,
            I => \N__44793\
        );

    \I__10336\ : LocalMux
    port map (
            O => \N__44802\,
            I => \N__44790\
        );

    \I__10335\ : LocalMux
    port map (
            O => \N__44799\,
            I => \N__44787\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__44796\,
            I => \N__44784\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__44793\,
            I => \N__44779\
        );

    \I__10332\ : Span12Mux_s6_v
    port map (
            O => \N__44790\,
            I => \N__44779\
        );

    \I__10331\ : Span4Mux_v
    port map (
            O => \N__44787\,
            I => \N__44774\
        );

    \I__10330\ : Span4Mux_h
    port map (
            O => \N__44784\,
            I => \N__44774\
        );

    \I__10329\ : Odrv12
    port map (
            O => \N__44779\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__10328\ : Odrv4
    port map (
            O => \N__44774\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__10327\ : InMux
    port map (
            O => \N__44769\,
            I => \N__44764\
        );

    \I__10326\ : InMux
    port map (
            O => \N__44768\,
            I => \N__44761\
        );

    \I__10325\ : InMux
    port map (
            O => \N__44767\,
            I => \N__44758\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__44764\,
            I => \N__44755\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__44761\,
            I => \N__44751\
        );

    \I__10322\ : LocalMux
    port map (
            O => \N__44758\,
            I => \N__44746\
        );

    \I__10321\ : Span4Mux_v
    port map (
            O => \N__44755\,
            I => \N__44746\
        );

    \I__10320\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44743\
        );

    \I__10319\ : Span4Mux_h
    port map (
            O => \N__44751\,
            I => \N__44740\
        );

    \I__10318\ : Sp12to4
    port map (
            O => \N__44746\,
            I => \N__44735\
        );

    \I__10317\ : LocalMux
    port map (
            O => \N__44743\,
            I => \N__44735\
        );

    \I__10316\ : Odrv4
    port map (
            O => \N__44740\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10315\ : Odrv12
    port map (
            O => \N__44735\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__10314\ : CascadeMux
    port map (
            O => \N__44730\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\
        );

    \I__10313\ : InMux
    port map (
            O => \N__44727\,
            I => \N__44724\
        );

    \I__10312\ : LocalMux
    port map (
            O => \N__44724\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__10311\ : InMux
    port map (
            O => \N__44721\,
            I => \N__44718\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__44718\,
            I => \N__44713\
        );

    \I__10309\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44710\
        );

    \I__10308\ : InMux
    port map (
            O => \N__44716\,
            I => \N__44707\
        );

    \I__10307\ : Span4Mux_v
    port map (
            O => \N__44713\,
            I => \N__44701\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__44710\,
            I => \N__44701\
        );

    \I__10305\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44698\
        );

    \I__10304\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44695\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__44701\,
            I => \N__44692\
        );

    \I__10302\ : Span4Mux_v
    port map (
            O => \N__44698\,
            I => \N__44689\
        );

    \I__10301\ : LocalMux
    port map (
            O => \N__44695\,
            I => \N__44686\
        );

    \I__10300\ : Span4Mux_h
    port map (
            O => \N__44692\,
            I => \N__44683\
        );

    \I__10299\ : Odrv4
    port map (
            O => \N__44689\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__10298\ : Odrv12
    port map (
            O => \N__44686\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__10297\ : Odrv4
    port map (
            O => \N__44683\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__10296\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44673\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__44673\,
            I => \N__44670\
        );

    \I__10294\ : Span4Mux_h
    port map (
            O => \N__44670\,
            I => \N__44667\
        );

    \I__10293\ : Odrv4
    port map (
            O => \N__44667\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__10292\ : CascadeMux
    port map (
            O => \N__44664\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__10291\ : CascadeMux
    port map (
            O => \N__44661\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__10290\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44655\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__44655\,
            I => \N__44652\
        );

    \I__10288\ : Odrv4
    port map (
            O => \N__44652\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\
        );

    \I__10287\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44646\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__44646\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__10285\ : InMux
    port map (
            O => \N__44643\,
            I => \N__44639\
        );

    \I__10284\ : InMux
    port map (
            O => \N__44642\,
            I => \N__44635\
        );

    \I__10283\ : LocalMux
    port map (
            O => \N__44639\,
            I => \N__44632\
        );

    \I__10282\ : InMux
    port map (
            O => \N__44638\,
            I => \N__44629\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__44635\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__44632\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__10279\ : LocalMux
    port map (
            O => \N__44629\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__10278\ : InMux
    port map (
            O => \N__44622\,
            I => \N__44618\
        );

    \I__10277\ : CascadeMux
    port map (
            O => \N__44621\,
            I => \N__44613\
        );

    \I__10276\ : LocalMux
    port map (
            O => \N__44618\,
            I => \N__44610\
        );

    \I__10275\ : InMux
    port map (
            O => \N__44617\,
            I => \N__44607\
        );

    \I__10274\ : InMux
    port map (
            O => \N__44616\,
            I => \N__44604\
        );

    \I__10273\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44601\
        );

    \I__10272\ : Span12Mux_h
    port map (
            O => \N__44610\,
            I => \N__44598\
        );

    \I__10271\ : LocalMux
    port map (
            O => \N__44607\,
            I => \N__44591\
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__44604\,
            I => \N__44591\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__44601\,
            I => \N__44591\
        );

    \I__10268\ : Odrv12
    port map (
            O => \N__44598\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10267\ : Odrv12
    port map (
            O => \N__44591\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__10266\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44583\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__44583\,
            I => \N__44580\
        );

    \I__10264\ : Span4Mux_h
    port map (
            O => \N__44580\,
            I => \N__44577\
        );

    \I__10263\ : Odrv4
    port map (
            O => \N__44577\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__10262\ : CascadeMux
    port map (
            O => \N__44574\,
            I => \N__44571\
        );

    \I__10261\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44567\
        );

    \I__10260\ : InMux
    port map (
            O => \N__44570\,
            I => \N__44564\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__44567\,
            I => \N__44558\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44558\
        );

    \I__10257\ : InMux
    port map (
            O => \N__44563\,
            I => \N__44555\
        );

    \I__10256\ : Span4Mux_h
    port map (
            O => \N__44558\,
            I => \N__44552\
        );

    \I__10255\ : LocalMux
    port map (
            O => \N__44555\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__44552\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__10253\ : InMux
    port map (
            O => \N__44547\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__10252\ : CascadeMux
    port map (
            O => \N__44544\,
            I => \N__44540\
        );

    \I__10251\ : CascadeMux
    port map (
            O => \N__44543\,
            I => \N__44537\
        );

    \I__10250\ : InMux
    port map (
            O => \N__44540\,
            I => \N__44531\
        );

    \I__10249\ : InMux
    port map (
            O => \N__44537\,
            I => \N__44531\
        );

    \I__10248\ : InMux
    port map (
            O => \N__44536\,
            I => \N__44528\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__44531\,
            I => \N__44525\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__44528\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10245\ : Odrv12
    port map (
            O => \N__44525\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__10244\ : InMux
    port map (
            O => \N__44520\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__10243\ : InMux
    port map (
            O => \N__44517\,
            I => \N__44513\
        );

    \I__10242\ : InMux
    port map (
            O => \N__44516\,
            I => \N__44510\
        );

    \I__10241\ : LocalMux
    port map (
            O => \N__44513\,
            I => \N__44507\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__44510\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10239\ : Odrv12
    port map (
            O => \N__44507\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__10238\ : InMux
    port map (
            O => \N__44502\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__10237\ : InMux
    port map (
            O => \N__44499\,
            I => \N__44463\
        );

    \I__10236\ : InMux
    port map (
            O => \N__44498\,
            I => \N__44463\
        );

    \I__10235\ : InMux
    port map (
            O => \N__44497\,
            I => \N__44463\
        );

    \I__10234\ : InMux
    port map (
            O => \N__44496\,
            I => \N__44454\
        );

    \I__10233\ : InMux
    port map (
            O => \N__44495\,
            I => \N__44454\
        );

    \I__10232\ : InMux
    port map (
            O => \N__44494\,
            I => \N__44454\
        );

    \I__10231\ : InMux
    port map (
            O => \N__44493\,
            I => \N__44454\
        );

    \I__10230\ : InMux
    port map (
            O => \N__44492\,
            I => \N__44445\
        );

    \I__10229\ : InMux
    port map (
            O => \N__44491\,
            I => \N__44445\
        );

    \I__10228\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44445\
        );

    \I__10227\ : InMux
    port map (
            O => \N__44489\,
            I => \N__44445\
        );

    \I__10226\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44436\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44436\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44486\,
            I => \N__44436\
        );

    \I__10223\ : InMux
    port map (
            O => \N__44485\,
            I => \N__44436\
        );

    \I__10222\ : InMux
    port map (
            O => \N__44484\,
            I => \N__44427\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44483\,
            I => \N__44427\
        );

    \I__10220\ : InMux
    port map (
            O => \N__44482\,
            I => \N__44427\
        );

    \I__10219\ : InMux
    port map (
            O => \N__44481\,
            I => \N__44427\
        );

    \I__10218\ : InMux
    port map (
            O => \N__44480\,
            I => \N__44420\
        );

    \I__10217\ : InMux
    port map (
            O => \N__44479\,
            I => \N__44420\
        );

    \I__10216\ : InMux
    port map (
            O => \N__44478\,
            I => \N__44420\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44411\
        );

    \I__10214\ : InMux
    port map (
            O => \N__44476\,
            I => \N__44411\
        );

    \I__10213\ : InMux
    port map (
            O => \N__44475\,
            I => \N__44411\
        );

    \I__10212\ : InMux
    port map (
            O => \N__44474\,
            I => \N__44411\
        );

    \I__10211\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44402\
        );

    \I__10210\ : InMux
    port map (
            O => \N__44472\,
            I => \N__44402\
        );

    \I__10209\ : InMux
    port map (
            O => \N__44471\,
            I => \N__44402\
        );

    \I__10208\ : InMux
    port map (
            O => \N__44470\,
            I => \N__44402\
        );

    \I__10207\ : LocalMux
    port map (
            O => \N__44463\,
            I => \N__44393\
        );

    \I__10206\ : LocalMux
    port map (
            O => \N__44454\,
            I => \N__44393\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__44445\,
            I => \N__44393\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__44436\,
            I => \N__44393\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__44427\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__44420\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10201\ : LocalMux
    port map (
            O => \N__44411\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44402\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10199\ : Odrv4
    port map (
            O => \N__44393\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44382\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__10197\ : InMux
    port map (
            O => \N__44379\,
            I => \N__44375\
        );

    \I__10196\ : InMux
    port map (
            O => \N__44378\,
            I => \N__44372\
        );

    \I__10195\ : LocalMux
    port map (
            O => \N__44375\,
            I => \N__44369\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__44372\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10193\ : Odrv12
    port map (
            O => \N__44369\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10192\ : CEMux
    port map (
            O => \N__44364\,
            I => \N__44360\
        );

    \I__10191\ : CEMux
    port map (
            O => \N__44363\,
            I => \N__44357\
        );

    \I__10190\ : LocalMux
    port map (
            O => \N__44360\,
            I => \N__44352\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__44357\,
            I => \N__44349\
        );

    \I__10188\ : CEMux
    port map (
            O => \N__44356\,
            I => \N__44346\
        );

    \I__10187\ : CEMux
    port map (
            O => \N__44355\,
            I => \N__44343\
        );

    \I__10186\ : Span4Mux_v
    port map (
            O => \N__44352\,
            I => \N__44338\
        );

    \I__10185\ : Span4Mux_v
    port map (
            O => \N__44349\,
            I => \N__44338\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__44346\,
            I => \N__44333\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__44343\,
            I => \N__44333\
        );

    \I__10182\ : Span4Mux_h
    port map (
            O => \N__44338\,
            I => \N__44328\
        );

    \I__10181\ : Span4Mux_v
    port map (
            O => \N__44333\,
            I => \N__44328\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__44328\,
            I => \current_shift_inst.timer_s1.N_163_i\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44322\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44317\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44314\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44311\
        );

    \I__10175\ : Span4Mux_v
    port map (
            O => \N__44317\,
            I => \N__44308\
        );

    \I__10174\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44305\
        );

    \I__10173\ : LocalMux
    port map (
            O => \N__44311\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__10172\ : Odrv4
    port map (
            O => \N__44308\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__10171\ : Odrv12
    port map (
            O => \N__44305\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44298\,
            I => \N__44293\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44297\,
            I => \N__44290\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44296\,
            I => \N__44287\
        );

    \I__10167\ : LocalMux
    port map (
            O => \N__44293\,
            I => \N__44283\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__44290\,
            I => \N__44278\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__44287\,
            I => \N__44278\
        );

    \I__10164\ : CascadeMux
    port map (
            O => \N__44286\,
            I => \N__44275\
        );

    \I__10163\ : Span4Mux_h
    port map (
            O => \N__44283\,
            I => \N__44272\
        );

    \I__10162\ : Span12Mux_h
    port map (
            O => \N__44278\,
            I => \N__44269\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44275\,
            I => \N__44266\
        );

    \I__10160\ : Odrv4
    port map (
            O => \N__44272\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10159\ : Odrv12
    port map (
            O => \N__44269\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44266\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__10157\ : InMux
    port map (
            O => \N__44259\,
            I => \N__44256\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44256\,
            I => \N__44252\
        );

    \I__10155\ : InMux
    port map (
            O => \N__44255\,
            I => \N__44248\
        );

    \I__10154\ : Span4Mux_h
    port map (
            O => \N__44252\,
            I => \N__44245\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44251\,
            I => \N__44242\
        );

    \I__10152\ : LocalMux
    port map (
            O => \N__44248\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10151\ : Odrv4
    port map (
            O => \N__44245\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10150\ : LocalMux
    port map (
            O => \N__44242\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__10149\ : InMux
    port map (
            O => \N__44235\,
            I => \N__44230\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44234\,
            I => \N__44227\
        );

    \I__10147\ : InMux
    port map (
            O => \N__44233\,
            I => \N__44224\
        );

    \I__10146\ : LocalMux
    port map (
            O => \N__44230\,
            I => \N__44221\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__44227\,
            I => \N__44218\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44224\,
            I => \N__44213\
        );

    \I__10143\ : Span4Mux_h
    port map (
            O => \N__44221\,
            I => \N__44213\
        );

    \I__10142\ : Span4Mux_h
    port map (
            O => \N__44218\,
            I => \N__44210\
        );

    \I__10141\ : Odrv4
    port map (
            O => \N__44213\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__10140\ : Odrv4
    port map (
            O => \N__44210\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__10139\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44202\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44202\,
            I => \N__44197\
        );

    \I__10137\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44194\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44200\,
            I => \N__44191\
        );

    \I__10135\ : Span4Mux_h
    port map (
            O => \N__44197\,
            I => \N__44188\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__44194\,
            I => \N__44185\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44191\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10132\ : Odrv4
    port map (
            O => \N__44188\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10131\ : Odrv12
    port map (
            O => \N__44185\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__10130\ : CascadeMux
    port map (
            O => \N__44178\,
            I => \N__44175\
        );

    \I__10129\ : InMux
    port map (
            O => \N__44175\,
            I => \N__44171\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44174\,
            I => \N__44168\
        );

    \I__10127\ : LocalMux
    port map (
            O => \N__44171\,
            I => \N__44162\
        );

    \I__10126\ : LocalMux
    port map (
            O => \N__44168\,
            I => \N__44162\
        );

    \I__10125\ : InMux
    port map (
            O => \N__44167\,
            I => \N__44159\
        );

    \I__10124\ : Span4Mux_h
    port map (
            O => \N__44162\,
            I => \N__44156\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__44159\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__10122\ : Odrv4
    port map (
            O => \N__44156\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44151\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__10120\ : CascadeMux
    port map (
            O => \N__44148\,
            I => \N__44144\
        );

    \I__10119\ : CascadeMux
    port map (
            O => \N__44147\,
            I => \N__44141\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44144\,
            I => \N__44135\
        );

    \I__10117\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44135\
        );

    \I__10116\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44132\
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44129\
        );

    \I__10114\ : LocalMux
    port map (
            O => \N__44132\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10113\ : Odrv12
    port map (
            O => \N__44129\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44124\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44121\,
            I => \N__44114\
        );

    \I__10110\ : InMux
    port map (
            O => \N__44120\,
            I => \N__44114\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44119\,
            I => \N__44111\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__44114\,
            I => \N__44108\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44111\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10106\ : Odrv12
    port map (
            O => \N__44108\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44103\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__10104\ : CascadeMux
    port map (
            O => \N__44100\,
            I => \N__44097\
        );

    \I__10103\ : InMux
    port map (
            O => \N__44097\,
            I => \N__44092\
        );

    \I__10102\ : InMux
    port map (
            O => \N__44096\,
            I => \N__44089\
        );

    \I__10101\ : InMux
    port map (
            O => \N__44095\,
            I => \N__44086\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__44092\,
            I => \N__44081\
        );

    \I__10099\ : LocalMux
    port map (
            O => \N__44089\,
            I => \N__44081\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44086\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10097\ : Odrv12
    port map (
            O => \N__44081\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__10096\ : InMux
    port map (
            O => \N__44076\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__10095\ : CascadeMux
    port map (
            O => \N__44073\,
            I => \N__44069\
        );

    \I__10094\ : CascadeMux
    port map (
            O => \N__44072\,
            I => \N__44066\
        );

    \I__10093\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44060\
        );

    \I__10092\ : InMux
    port map (
            O => \N__44066\,
            I => \N__44060\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44065\,
            I => \N__44057\
        );

    \I__10090\ : LocalMux
    port map (
            O => \N__44060\,
            I => \N__44054\
        );

    \I__10089\ : LocalMux
    port map (
            O => \N__44057\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10088\ : Odrv12
    port map (
            O => \N__44054\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__10087\ : InMux
    port map (
            O => \N__44049\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__10086\ : InMux
    port map (
            O => \N__44046\,
            I => \N__44039\
        );

    \I__10085\ : InMux
    port map (
            O => \N__44045\,
            I => \N__44039\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44044\,
            I => \N__44036\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44039\,
            I => \N__44033\
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__44036\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__10081\ : Odrv12
    port map (
            O => \N__44033\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__10080\ : InMux
    port map (
            O => \N__44028\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__10079\ : CascadeMux
    port map (
            O => \N__44025\,
            I => \N__44022\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44022\,
            I => \N__44018\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44021\,
            I => \N__44015\
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__44018\,
            I => \N__44009\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44015\,
            I => \N__44009\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44014\,
            I => \N__44006\
        );

    \I__10073\ : Span4Mux_v
    port map (
            O => \N__44009\,
            I => \N__44003\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__44006\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__44003\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__10070\ : InMux
    port map (
            O => \N__43998\,
            I => \bfn_17_22_0_\
        );

    \I__10069\ : InMux
    port map (
            O => \N__43995\,
            I => \N__43991\
        );

    \I__10068\ : CascadeMux
    port map (
            O => \N__43994\,
            I => \N__43988\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__43991\,
            I => \N__43984\
        );

    \I__10066\ : InMux
    port map (
            O => \N__43988\,
            I => \N__43981\
        );

    \I__10065\ : InMux
    port map (
            O => \N__43987\,
            I => \N__43978\
        );

    \I__10064\ : Span4Mux_h
    port map (
            O => \N__43984\,
            I => \N__43975\
        );

    \I__10063\ : LocalMux
    port map (
            O => \N__43981\,
            I => \N__43972\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__43978\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10061\ : Odrv4
    port map (
            O => \N__43975\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10060\ : Odrv12
    port map (
            O => \N__43972\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__10059\ : InMux
    port map (
            O => \N__43965\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__10058\ : CascadeMux
    port map (
            O => \N__43962\,
            I => \N__43959\
        );

    \I__10057\ : InMux
    port map (
            O => \N__43959\,
            I => \N__43956\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__43956\,
            I => \N__43951\
        );

    \I__10055\ : InMux
    port map (
            O => \N__43955\,
            I => \N__43948\
        );

    \I__10054\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43945\
        );

    \I__10053\ : Span4Mux_h
    port map (
            O => \N__43951\,
            I => \N__43942\
        );

    \I__10052\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43939\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__43945\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10050\ : Odrv4
    port map (
            O => \N__43942\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10049\ : Odrv12
    port map (
            O => \N__43939\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__10048\ : InMux
    port map (
            O => \N__43932\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__10047\ : InMux
    port map (
            O => \N__43929\,
            I => \N__43922\
        );

    \I__10046\ : InMux
    port map (
            O => \N__43928\,
            I => \N__43922\
        );

    \I__10045\ : InMux
    port map (
            O => \N__43927\,
            I => \N__43919\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__43922\,
            I => \N__43916\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__43919\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__10042\ : Odrv12
    port map (
            O => \N__43916\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__10041\ : InMux
    port map (
            O => \N__43911\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__10040\ : InMux
    port map (
            O => \N__43908\,
            I => \N__43902\
        );

    \I__10039\ : InMux
    port map (
            O => \N__43907\,
            I => \N__43902\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__43902\,
            I => \N__43898\
        );

    \I__10037\ : InMux
    port map (
            O => \N__43901\,
            I => \N__43895\
        );

    \I__10036\ : Span4Mux_h
    port map (
            O => \N__43898\,
            I => \N__43892\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__43895\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10034\ : Odrv4
    port map (
            O => \N__43892\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__10033\ : InMux
    port map (
            O => \N__43887\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__10032\ : CascadeMux
    port map (
            O => \N__43884\,
            I => \N__43880\
        );

    \I__10031\ : InMux
    port map (
            O => \N__43883\,
            I => \N__43876\
        );

    \I__10030\ : InMux
    port map (
            O => \N__43880\,
            I => \N__43873\
        );

    \I__10029\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43870\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__43876\,
            I => \N__43865\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__43873\,
            I => \N__43865\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__43870\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10025\ : Odrv12
    port map (
            O => \N__43865\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__10024\ : InMux
    port map (
            O => \N__43860\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__10023\ : CascadeMux
    port map (
            O => \N__43857\,
            I => \N__43853\
        );

    \I__10022\ : CascadeMux
    port map (
            O => \N__43856\,
            I => \N__43850\
        );

    \I__10021\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43845\
        );

    \I__10020\ : InMux
    port map (
            O => \N__43850\,
            I => \N__43845\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__43845\,
            I => \N__43841\
        );

    \I__10018\ : InMux
    port map (
            O => \N__43844\,
            I => \N__43838\
        );

    \I__10017\ : Span4Mux_h
    port map (
            O => \N__43841\,
            I => \N__43835\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__43838\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10015\ : Odrv4
    port map (
            O => \N__43835\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__10014\ : InMux
    port map (
            O => \N__43830\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__10013\ : CascadeMux
    port map (
            O => \N__43827\,
            I => \N__43823\
        );

    \I__10012\ : CascadeMux
    port map (
            O => \N__43826\,
            I => \N__43820\
        );

    \I__10011\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43815\
        );

    \I__10010\ : InMux
    port map (
            O => \N__43820\,
            I => \N__43815\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__43815\,
            I => \N__43811\
        );

    \I__10008\ : InMux
    port map (
            O => \N__43814\,
            I => \N__43808\
        );

    \I__10007\ : Span4Mux_v
    port map (
            O => \N__43811\,
            I => \N__43805\
        );

    \I__10006\ : LocalMux
    port map (
            O => \N__43808\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10005\ : Odrv4
    port map (
            O => \N__43805\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__10004\ : InMux
    port map (
            O => \N__43800\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__10003\ : InMux
    port map (
            O => \N__43797\,
            I => \N__43791\
        );

    \I__10002\ : InMux
    port map (
            O => \N__43796\,
            I => \N__43791\
        );

    \I__10001\ : LocalMux
    port map (
            O => \N__43791\,
            I => \N__43787\
        );

    \I__10000\ : InMux
    port map (
            O => \N__43790\,
            I => \N__43784\
        );

    \I__9999\ : Span4Mux_v
    port map (
            O => \N__43787\,
            I => \N__43781\
        );

    \I__9998\ : LocalMux
    port map (
            O => \N__43784\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9997\ : Odrv4
    port map (
            O => \N__43781\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9996\ : InMux
    port map (
            O => \N__43776\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__9995\ : CascadeMux
    port map (
            O => \N__43773\,
            I => \N__43770\
        );

    \I__9994\ : InMux
    port map (
            O => \N__43770\,
            I => \N__43766\
        );

    \I__9993\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43763\
        );

    \I__9992\ : LocalMux
    port map (
            O => \N__43766\,
            I => \N__43757\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__43763\,
            I => \N__43757\
        );

    \I__9990\ : InMux
    port map (
            O => \N__43762\,
            I => \N__43754\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__43757\,
            I => \N__43751\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__43754\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9987\ : Odrv4
    port map (
            O => \N__43751\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9986\ : InMux
    port map (
            O => \N__43746\,
            I => \bfn_17_21_0_\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__43743\,
            I => \N__43739\
        );

    \I__9984\ : InMux
    port map (
            O => \N__43742\,
            I => \N__43736\
        );

    \I__9983\ : InMux
    port map (
            O => \N__43739\,
            I => \N__43733\
        );

    \I__9982\ : LocalMux
    port map (
            O => \N__43736\,
            I => \N__43729\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__43733\,
            I => \N__43726\
        );

    \I__9980\ : InMux
    port map (
            O => \N__43732\,
            I => \N__43723\
        );

    \I__9979\ : Span4Mux_v
    port map (
            O => \N__43729\,
            I => \N__43718\
        );

    \I__9978\ : Span4Mux_v
    port map (
            O => \N__43726\,
            I => \N__43718\
        );

    \I__9977\ : LocalMux
    port map (
            O => \N__43723\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9976\ : Odrv4
    port map (
            O => \N__43718\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9975\ : InMux
    port map (
            O => \N__43713\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__9974\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43707\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__43707\,
            I => \N__43703\
        );

    \I__9972\ : InMux
    port map (
            O => \N__43706\,
            I => \N__43699\
        );

    \I__9971\ : Span4Mux_h
    port map (
            O => \N__43703\,
            I => \N__43696\
        );

    \I__9970\ : InMux
    port map (
            O => \N__43702\,
            I => \N__43693\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__43699\,
            I => \N__43690\
        );

    \I__9968\ : Odrv4
    port map (
            O => \N__43696\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__43693\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9966\ : Odrv12
    port map (
            O => \N__43690\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__9965\ : InMux
    port map (
            O => \N__43683\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__9964\ : InMux
    port map (
            O => \N__43680\,
            I => \N__43676\
        );

    \I__9963\ : CascadeMux
    port map (
            O => \N__43679\,
            I => \N__43673\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__43676\,
            I => \N__43669\
        );

    \I__9961\ : InMux
    port map (
            O => \N__43673\,
            I => \N__43666\
        );

    \I__9960\ : InMux
    port map (
            O => \N__43672\,
            I => \N__43663\
        );

    \I__9959\ : Sp12to4
    port map (
            O => \N__43669\,
            I => \N__43658\
        );

    \I__9958\ : LocalMux
    port map (
            O => \N__43666\,
            I => \N__43658\
        );

    \I__9957\ : LocalMux
    port map (
            O => \N__43663\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9956\ : Odrv12
    port map (
            O => \N__43658\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9955\ : InMux
    port map (
            O => \N__43653\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__9954\ : CascadeMux
    port map (
            O => \N__43650\,
            I => \N__43646\
        );

    \I__9953\ : InMux
    port map (
            O => \N__43649\,
            I => \N__43643\
        );

    \I__9952\ : InMux
    port map (
            O => \N__43646\,
            I => \N__43640\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__43643\,
            I => \N__43634\
        );

    \I__9950\ : LocalMux
    port map (
            O => \N__43640\,
            I => \N__43634\
        );

    \I__9949\ : InMux
    port map (
            O => \N__43639\,
            I => \N__43631\
        );

    \I__9948\ : Span4Mux_v
    port map (
            O => \N__43634\,
            I => \N__43628\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__43631\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9946\ : Odrv4
    port map (
            O => \N__43628\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9945\ : InMux
    port map (
            O => \N__43623\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__9944\ : CascadeMux
    port map (
            O => \N__43620\,
            I => \N__43616\
        );

    \I__9943\ : CascadeMux
    port map (
            O => \N__43619\,
            I => \N__43613\
        );

    \I__9942\ : InMux
    port map (
            O => \N__43616\,
            I => \N__43608\
        );

    \I__9941\ : InMux
    port map (
            O => \N__43613\,
            I => \N__43608\
        );

    \I__9940\ : LocalMux
    port map (
            O => \N__43608\,
            I => \N__43604\
        );

    \I__9939\ : InMux
    port map (
            O => \N__43607\,
            I => \N__43601\
        );

    \I__9938\ : Span4Mux_v
    port map (
            O => \N__43604\,
            I => \N__43598\
        );

    \I__9937\ : LocalMux
    port map (
            O => \N__43601\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9936\ : Odrv4
    port map (
            O => \N__43598\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9935\ : InMux
    port map (
            O => \N__43593\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__9934\ : CascadeMux
    port map (
            O => \N__43590\,
            I => \N__43586\
        );

    \I__9933\ : CascadeMux
    port map (
            O => \N__43589\,
            I => \N__43583\
        );

    \I__9932\ : InMux
    port map (
            O => \N__43586\,
            I => \N__43578\
        );

    \I__9931\ : InMux
    port map (
            O => \N__43583\,
            I => \N__43578\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__43578\,
            I => \N__43574\
        );

    \I__9929\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43571\
        );

    \I__9928\ : Span4Mux_h
    port map (
            O => \N__43574\,
            I => \N__43568\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__43571\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9926\ : Odrv4
    port map (
            O => \N__43568\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9925\ : InMux
    port map (
            O => \N__43563\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__9924\ : InMux
    port map (
            O => \N__43560\,
            I => \N__43554\
        );

    \I__9923\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43554\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__43554\,
            I => \N__43550\
        );

    \I__9921\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43547\
        );

    \I__9920\ : Span4Mux_v
    port map (
            O => \N__43550\,
            I => \N__43544\
        );

    \I__9919\ : LocalMux
    port map (
            O => \N__43547\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9918\ : Odrv4
    port map (
            O => \N__43544\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9917\ : InMux
    port map (
            O => \N__43539\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__9916\ : CascadeMux
    port map (
            O => \N__43536\,
            I => \N__43533\
        );

    \I__9915\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43529\
        );

    \I__9914\ : InMux
    port map (
            O => \N__43532\,
            I => \N__43526\
        );

    \I__9913\ : LocalMux
    port map (
            O => \N__43529\,
            I => \N__43520\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__43526\,
            I => \N__43520\
        );

    \I__9911\ : InMux
    port map (
            O => \N__43525\,
            I => \N__43517\
        );

    \I__9910\ : Span4Mux_v
    port map (
            O => \N__43520\,
            I => \N__43514\
        );

    \I__9909\ : LocalMux
    port map (
            O => \N__43517\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9908\ : Odrv4
    port map (
            O => \N__43514\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9907\ : InMux
    port map (
            O => \N__43509\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__9906\ : CascadeMux
    port map (
            O => \N__43506\,
            I => \N__43502\
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__43505\,
            I => \N__43499\
        );

    \I__9904\ : InMux
    port map (
            O => \N__43502\,
            I => \N__43496\
        );

    \I__9903\ : InMux
    port map (
            O => \N__43499\,
            I => \N__43493\
        );

    \I__9902\ : LocalMux
    port map (
            O => \N__43496\,
            I => \N__43487\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43493\,
            I => \N__43487\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43484\
        );

    \I__9899\ : Span4Mux_v
    port map (
            O => \N__43487\,
            I => \N__43481\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43484\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__43481\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9896\ : InMux
    port map (
            O => \N__43476\,
            I => \bfn_17_20_0_\
        );

    \I__9895\ : InMux
    port map (
            O => \N__43473\,
            I => \N__43468\
        );

    \I__9894\ : InMux
    port map (
            O => \N__43472\,
            I => \N__43465\
        );

    \I__9893\ : InMux
    port map (
            O => \N__43471\,
            I => \N__43462\
        );

    \I__9892\ : LocalMux
    port map (
            O => \N__43468\,
            I => \N__43459\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__43465\,
            I => \N__43456\
        );

    \I__9890\ : LocalMux
    port map (
            O => \N__43462\,
            I => \N__43453\
        );

    \I__9889\ : Span4Mux_h
    port map (
            O => \N__43459\,
            I => \N__43449\
        );

    \I__9888\ : Span4Mux_h
    port map (
            O => \N__43456\,
            I => \N__43446\
        );

    \I__9887\ : Span4Mux_h
    port map (
            O => \N__43453\,
            I => \N__43443\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43452\,
            I => \N__43440\
        );

    \I__9885\ : Odrv4
    port map (
            O => \N__43449\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9884\ : Odrv4
    port map (
            O => \N__43446\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9883\ : Odrv4
    port map (
            O => \N__43443\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43440\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9881\ : InMux
    port map (
            O => \N__43431\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__9880\ : InMux
    port map (
            O => \N__43428\,
            I => \N__43423\
        );

    \I__9879\ : InMux
    port map (
            O => \N__43427\,
            I => \N__43420\
        );

    \I__9878\ : InMux
    port map (
            O => \N__43426\,
            I => \N__43417\
        );

    \I__9877\ : LocalMux
    port map (
            O => \N__43423\,
            I => \N__43413\
        );

    \I__9876\ : LocalMux
    port map (
            O => \N__43420\,
            I => \N__43408\
        );

    \I__9875\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43408\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43416\,
            I => \N__43405\
        );

    \I__9873\ : Span4Mux_v
    port map (
            O => \N__43413\,
            I => \N__43398\
        );

    \I__9872\ : Span4Mux_v
    port map (
            O => \N__43408\,
            I => \N__43398\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43405\,
            I => \N__43398\
        );

    \I__9870\ : Odrv4
    port map (
            O => \N__43398\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9869\ : InMux
    port map (
            O => \N__43395\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__9868\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43387\
        );

    \I__9867\ : InMux
    port map (
            O => \N__43391\,
            I => \N__43384\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43390\,
            I => \N__43381\
        );

    \I__9865\ : LocalMux
    port map (
            O => \N__43387\,
            I => \N__43376\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__43384\,
            I => \N__43376\
        );

    \I__9863\ : LocalMux
    port map (
            O => \N__43381\,
            I => \N__43373\
        );

    \I__9862\ : Span4Mux_v
    port map (
            O => \N__43376\,
            I => \N__43369\
        );

    \I__9861\ : Span4Mux_h
    port map (
            O => \N__43373\,
            I => \N__43366\
        );

    \I__9860\ : InMux
    port map (
            O => \N__43372\,
            I => \N__43363\
        );

    \I__9859\ : Odrv4
    port map (
            O => \N__43369\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9858\ : Odrv4
    port map (
            O => \N__43366\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43363\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9856\ : InMux
    port map (
            O => \N__43356\,
            I => \bfn_17_18_0_\
        );

    \I__9855\ : InMux
    port map (
            O => \N__43353\,
            I => \N__43347\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43352\,
            I => \N__43347\
        );

    \I__9853\ : LocalMux
    port map (
            O => \N__43347\,
            I => \N__43343\
        );

    \I__9852\ : InMux
    port map (
            O => \N__43346\,
            I => \N__43340\
        );

    \I__9851\ : Span4Mux_v
    port map (
            O => \N__43343\,
            I => \N__43335\
        );

    \I__9850\ : LocalMux
    port map (
            O => \N__43340\,
            I => \N__43335\
        );

    \I__9849\ : Span4Mux_h
    port map (
            O => \N__43335\,
            I => \N__43331\
        );

    \I__9848\ : InMux
    port map (
            O => \N__43334\,
            I => \N__43328\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__43331\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9846\ : LocalMux
    port map (
            O => \N__43328\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43323\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43320\,
            I => \N__43316\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43319\,
            I => \N__43313\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__43316\,
            I => \N__43307\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43313\,
            I => \N__43307\
        );

    \I__9840\ : InMux
    port map (
            O => \N__43312\,
            I => \N__43304\
        );

    \I__9839\ : Span4Mux_v
    port map (
            O => \N__43307\,
            I => \N__43298\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43304\,
            I => \N__43298\
        );

    \I__9837\ : InMux
    port map (
            O => \N__43303\,
            I => \N__43295\
        );

    \I__9836\ : Span4Mux_h
    port map (
            O => \N__43298\,
            I => \N__43292\
        );

    \I__9835\ : LocalMux
    port map (
            O => \N__43295\,
            I => \N__43289\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__43292\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9833\ : Odrv12
    port map (
            O => \N__43289\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43284\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__9831\ : InMux
    port map (
            O => \N__43281\,
            I => \N__43277\
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__43280\,
            I => \N__43274\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__43277\,
            I => \N__43270\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43267\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43264\
        );

    \I__9826\ : Span4Mux_v
    port map (
            O => \N__43270\,
            I => \N__43261\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__43267\,
            I => \N__43258\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__43264\,
            I => \N__43255\
        );

    \I__9823\ : Span4Mux_h
    port map (
            O => \N__43261\,
            I => \N__43249\
        );

    \I__9822\ : Span4Mux_v
    port map (
            O => \N__43258\,
            I => \N__43249\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__43255\,
            I => \N__43246\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43254\,
            I => \N__43243\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__43249\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9818\ : Odrv4
    port map (
            O => \N__43246\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__43243\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43236\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__9815\ : CEMux
    port map (
            O => \N__43233\,
            I => \N__43209\
        );

    \I__9814\ : CEMux
    port map (
            O => \N__43232\,
            I => \N__43209\
        );

    \I__9813\ : CEMux
    port map (
            O => \N__43231\,
            I => \N__43209\
        );

    \I__9812\ : CEMux
    port map (
            O => \N__43230\,
            I => \N__43209\
        );

    \I__9811\ : CEMux
    port map (
            O => \N__43229\,
            I => \N__43209\
        );

    \I__9810\ : CEMux
    port map (
            O => \N__43228\,
            I => \N__43209\
        );

    \I__9809\ : CEMux
    port map (
            O => \N__43227\,
            I => \N__43209\
        );

    \I__9808\ : CEMux
    port map (
            O => \N__43226\,
            I => \N__43209\
        );

    \I__9807\ : GlobalMux
    port map (
            O => \N__43209\,
            I => \N__43206\
        );

    \I__9806\ : gio2CtrlBuf
    port map (
            O => \N__43206\,
            I => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \I__9805\ : InMux
    port map (
            O => \N__43203\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43200\,
            I => \N__43197\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43197\,
            I => \N__43194\
        );

    \I__9802\ : Span4Mux_v
    port map (
            O => \N__43194\,
            I => \N__43189\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43193\,
            I => \N__43186\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43192\,
            I => \N__43183\
        );

    \I__9799\ : Span4Mux_v
    port map (
            O => \N__43189\,
            I => \N__43176\
        );

    \I__9798\ : LocalMux
    port map (
            O => \N__43186\,
            I => \N__43176\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__43183\,
            I => \N__43176\
        );

    \I__9796\ : Span4Mux_v
    port map (
            O => \N__43176\,
            I => \N__43173\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__43173\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__9794\ : InMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__9793\ : LocalMux
    port map (
            O => \N__43167\,
            I => \N__43163\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43166\,
            I => \N__43159\
        );

    \I__9791\ : Span12Mux_v
    port map (
            O => \N__43163\,
            I => \N__43156\
        );

    \I__9790\ : InMux
    port map (
            O => \N__43162\,
            I => \N__43153\
        );

    \I__9789\ : LocalMux
    port map (
            O => \N__43159\,
            I => \N__43150\
        );

    \I__9788\ : Odrv12
    port map (
            O => \N__43156\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43153\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9786\ : Odrv12
    port map (
            O => \N__43150\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43143\,
            I => \bfn_17_19_0_\
        );

    \I__9784\ : CascadeMux
    port map (
            O => \N__43140\,
            I => \N__43136\
        );

    \I__9783\ : InMux
    port map (
            O => \N__43139\,
            I => \N__43133\
        );

    \I__9782\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43129\
        );

    \I__9781\ : LocalMux
    port map (
            O => \N__43133\,
            I => \N__43126\
        );

    \I__9780\ : InMux
    port map (
            O => \N__43132\,
            I => \N__43123\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__43129\,
            I => \N__43120\
        );

    \I__9778\ : Span4Mux_h
    port map (
            O => \N__43126\,
            I => \N__43115\
        );

    \I__9777\ : LocalMux
    port map (
            O => \N__43123\,
            I => \N__43115\
        );

    \I__9776\ : Span4Mux_h
    port map (
            O => \N__43120\,
            I => \N__43111\
        );

    \I__9775\ : Span4Mux_v
    port map (
            O => \N__43115\,
            I => \N__43108\
        );

    \I__9774\ : InMux
    port map (
            O => \N__43114\,
            I => \N__43105\
        );

    \I__9773\ : Odrv4
    port map (
            O => \N__43111\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9772\ : Odrv4
    port map (
            O => \N__43108\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9771\ : LocalMux
    port map (
            O => \N__43105\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9770\ : InMux
    port map (
            O => \N__43098\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__9769\ : CascadeMux
    port map (
            O => \N__43095\,
            I => \N__43092\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43092\,
            I => \N__43089\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43089\,
            I => \N__43084\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43081\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43087\,
            I => \N__43078\
        );

    \I__9764\ : Span4Mux_v
    port map (
            O => \N__43084\,
            I => \N__43075\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43081\,
            I => \N__43070\
        );

    \I__9762\ : LocalMux
    port map (
            O => \N__43078\,
            I => \N__43070\
        );

    \I__9761\ : Span4Mux_h
    port map (
            O => \N__43075\,
            I => \N__43066\
        );

    \I__9760\ : Span4Mux_h
    port map (
            O => \N__43070\,
            I => \N__43063\
        );

    \I__9759\ : InMux
    port map (
            O => \N__43069\,
            I => \N__43060\
        );

    \I__9758\ : Odrv4
    port map (
            O => \N__43066\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9757\ : Odrv4
    port map (
            O => \N__43063\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43060\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9755\ : InMux
    port map (
            O => \N__43053\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__9754\ : CascadeMux
    port map (
            O => \N__43050\,
            I => \N__43047\
        );

    \I__9753\ : InMux
    port map (
            O => \N__43047\,
            I => \N__43043\
        );

    \I__9752\ : InMux
    port map (
            O => \N__43046\,
            I => \N__43039\
        );

    \I__9751\ : LocalMux
    port map (
            O => \N__43043\,
            I => \N__43036\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43042\,
            I => \N__43033\
        );

    \I__9749\ : LocalMux
    port map (
            O => \N__43039\,
            I => \N__43030\
        );

    \I__9748\ : Span4Mux_v
    port map (
            O => \N__43036\,
            I => \N__43024\
        );

    \I__9747\ : LocalMux
    port map (
            O => \N__43033\,
            I => \N__43024\
        );

    \I__9746\ : Span4Mux_h
    port map (
            O => \N__43030\,
            I => \N__43021\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43029\,
            I => \N__43018\
        );

    \I__9744\ : Odrv4
    port map (
            O => \N__43024\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__9743\ : Odrv4
    port map (
            O => \N__43021\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43018\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__9741\ : InMux
    port map (
            O => \N__43011\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__9740\ : CascadeMux
    port map (
            O => \N__43008\,
            I => \N__43004\
        );

    \I__9739\ : InMux
    port map (
            O => \N__43007\,
            I => \N__43001\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43004\,
            I => \N__42998\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__43001\,
            I => \N__42994\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__42998\,
            I => \N__42991\
        );

    \I__9735\ : InMux
    port map (
            O => \N__42997\,
            I => \N__42988\
        );

    \I__9734\ : Span4Mux_h
    port map (
            O => \N__42994\,
            I => \N__42981\
        );

    \I__9733\ : Span4Mux_v
    port map (
            O => \N__42991\,
            I => \N__42981\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__42988\,
            I => \N__42981\
        );

    \I__9731\ : Span4Mux_h
    port map (
            O => \N__42981\,
            I => \N__42977\
        );

    \I__9730\ : InMux
    port map (
            O => \N__42980\,
            I => \N__42974\
        );

    \I__9729\ : Odrv4
    port map (
            O => \N__42977\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__42974\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9727\ : InMux
    port map (
            O => \N__42969\,
            I => \bfn_17_17_0_\
        );

    \I__9726\ : InMux
    port map (
            O => \N__42966\,
            I => \N__42960\
        );

    \I__9725\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42960\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__42960\,
            I => \N__42956\
        );

    \I__9723\ : InMux
    port map (
            O => \N__42959\,
            I => \N__42953\
        );

    \I__9722\ : Span4Mux_v
    port map (
            O => \N__42956\,
            I => \N__42948\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__42953\,
            I => \N__42948\
        );

    \I__9720\ : Span4Mux_h
    port map (
            O => \N__42948\,
            I => \N__42944\
        );

    \I__9719\ : InMux
    port map (
            O => \N__42947\,
            I => \N__42941\
        );

    \I__9718\ : Odrv4
    port map (
            O => \N__42944\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__42941\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9716\ : InMux
    port map (
            O => \N__42936\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__9715\ : InMux
    port map (
            O => \N__42933\,
            I => \N__42928\
        );

    \I__9714\ : InMux
    port map (
            O => \N__42932\,
            I => \N__42925\
        );

    \I__9713\ : InMux
    port map (
            O => \N__42931\,
            I => \N__42922\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__42928\,
            I => \N__42917\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__42925\,
            I => \N__42917\
        );

    \I__9710\ : LocalMux
    port map (
            O => \N__42922\,
            I => \N__42914\
        );

    \I__9709\ : Span4Mux_h
    port map (
            O => \N__42917\,
            I => \N__42910\
        );

    \I__9708\ : Span4Mux_h
    port map (
            O => \N__42914\,
            I => \N__42907\
        );

    \I__9707\ : InMux
    port map (
            O => \N__42913\,
            I => \N__42904\
        );

    \I__9706\ : Odrv4
    port map (
            O => \N__42910\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__42907\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9704\ : LocalMux
    port map (
            O => \N__42904\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__9703\ : InMux
    port map (
            O => \N__42897\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__9702\ : InMux
    port map (
            O => \N__42894\,
            I => \N__42889\
        );

    \I__9701\ : InMux
    port map (
            O => \N__42893\,
            I => \N__42886\
        );

    \I__9700\ : InMux
    port map (
            O => \N__42892\,
            I => \N__42883\
        );

    \I__9699\ : LocalMux
    port map (
            O => \N__42889\,
            I => \N__42880\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__42886\,
            I => \N__42875\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__42883\,
            I => \N__42875\
        );

    \I__9696\ : Span4Mux_v
    port map (
            O => \N__42880\,
            I => \N__42869\
        );

    \I__9695\ : Span4Mux_v
    port map (
            O => \N__42875\,
            I => \N__42869\
        );

    \I__9694\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42866\
        );

    \I__9693\ : Odrv4
    port map (
            O => \N__42869\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9692\ : LocalMux
    port map (
            O => \N__42866\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__9691\ : InMux
    port map (
            O => \N__42861\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__9690\ : InMux
    port map (
            O => \N__42858\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__9689\ : InMux
    port map (
            O => \N__42855\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__9688\ : CascadeMux
    port map (
            O => \N__42852\,
            I => \N__42848\
        );

    \I__9687\ : CascadeMux
    port map (
            O => \N__42851\,
            I => \N__42845\
        );

    \I__9686\ : InMux
    port map (
            O => \N__42848\,
            I => \N__42842\
        );

    \I__9685\ : InMux
    port map (
            O => \N__42845\,
            I => \N__42839\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__42842\,
            I => \N__42835\
        );

    \I__9683\ : LocalMux
    port map (
            O => \N__42839\,
            I => \N__42832\
        );

    \I__9682\ : InMux
    port map (
            O => \N__42838\,
            I => \N__42829\
        );

    \I__9681\ : Span4Mux_v
    port map (
            O => \N__42835\,
            I => \N__42826\
        );

    \I__9680\ : Span4Mux_v
    port map (
            O => \N__42832\,
            I => \N__42821\
        );

    \I__9679\ : LocalMux
    port map (
            O => \N__42829\,
            I => \N__42821\
        );

    \I__9678\ : Span4Mux_h
    port map (
            O => \N__42826\,
            I => \N__42817\
        );

    \I__9677\ : Span4Mux_h
    port map (
            O => \N__42821\,
            I => \N__42814\
        );

    \I__9676\ : InMux
    port map (
            O => \N__42820\,
            I => \N__42811\
        );

    \I__9675\ : Odrv4
    port map (
            O => \N__42817\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9674\ : Odrv4
    port map (
            O => \N__42814\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__42811\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__9672\ : InMux
    port map (
            O => \N__42804\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__9671\ : CascadeMux
    port map (
            O => \N__42801\,
            I => \N__42797\
        );

    \I__9670\ : InMux
    port map (
            O => \N__42800\,
            I => \N__42793\
        );

    \I__9669\ : InMux
    port map (
            O => \N__42797\,
            I => \N__42790\
        );

    \I__9668\ : InMux
    port map (
            O => \N__42796\,
            I => \N__42787\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__42793\,
            I => \N__42784\
        );

    \I__9666\ : LocalMux
    port map (
            O => \N__42790\,
            I => \N__42781\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__42787\,
            I => \N__42778\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__42784\,
            I => \N__42774\
        );

    \I__9663\ : Span4Mux_v
    port map (
            O => \N__42781\,
            I => \N__42769\
        );

    \I__9662\ : Span4Mux_v
    port map (
            O => \N__42778\,
            I => \N__42769\
        );

    \I__9661\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42766\
        );

    \I__9660\ : Odrv4
    port map (
            O => \N__42774\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9659\ : Odrv4
    port map (
            O => \N__42769\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__42766\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9657\ : InMux
    port map (
            O => \N__42759\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__9656\ : CascadeMux
    port map (
            O => \N__42756\,
            I => \N__42752\
        );

    \I__9655\ : InMux
    port map (
            O => \N__42755\,
            I => \N__42749\
        );

    \I__9654\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42746\
        );

    \I__9653\ : LocalMux
    port map (
            O => \N__42749\,
            I => \N__42743\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__42746\,
            I => \N__42739\
        );

    \I__9651\ : Span4Mux_v
    port map (
            O => \N__42743\,
            I => \N__42736\
        );

    \I__9650\ : InMux
    port map (
            O => \N__42742\,
            I => \N__42733\
        );

    \I__9649\ : Span4Mux_v
    port map (
            O => \N__42739\,
            I => \N__42725\
        );

    \I__9648\ : Span4Mux_h
    port map (
            O => \N__42736\,
            I => \N__42725\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__42733\,
            I => \N__42725\
        );

    \I__9646\ : InMux
    port map (
            O => \N__42732\,
            I => \N__42722\
        );

    \I__9645\ : Odrv4
    port map (
            O => \N__42725\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9644\ : LocalMux
    port map (
            O => \N__42722\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__9643\ : InMux
    port map (
            O => \N__42717\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__9642\ : CascadeMux
    port map (
            O => \N__42714\,
            I => \N__42711\
        );

    \I__9641\ : InMux
    port map (
            O => \N__42711\,
            I => \N__42706\
        );

    \I__9640\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42701\
        );

    \I__9639\ : InMux
    port map (
            O => \N__42709\,
            I => \N__42701\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__42706\,
            I => \N__42698\
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__42701\,
            I => \N__42695\
        );

    \I__9636\ : Span12Mux_v
    port map (
            O => \N__42698\,
            I => \N__42691\
        );

    \I__9635\ : Span4Mux_v
    port map (
            O => \N__42695\,
            I => \N__42688\
        );

    \I__9634\ : InMux
    port map (
            O => \N__42694\,
            I => \N__42685\
        );

    \I__9633\ : Odrv12
    port map (
            O => \N__42691\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__9632\ : Odrv4
    port map (
            O => \N__42688\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__42685\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__9630\ : InMux
    port map (
            O => \N__42678\,
            I => \bfn_17_16_0_\
        );

    \I__9629\ : InMux
    port map (
            O => \N__42675\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__42672\,
            I => \N__42667\
        );

    \I__9627\ : InMux
    port map (
            O => \N__42671\,
            I => \N__42664\
        );

    \I__9626\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42661\
        );

    \I__9625\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42658\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__42664\,
            I => \N__42655\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__42661\,
            I => \N__42652\
        );

    \I__9622\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42648\
        );

    \I__9621\ : Span4Mux_v
    port map (
            O => \N__42655\,
            I => \N__42643\
        );

    \I__9620\ : Span4Mux_v
    port map (
            O => \N__42652\,
            I => \N__42643\
        );

    \I__9619\ : InMux
    port map (
            O => \N__42651\,
            I => \N__42640\
        );

    \I__9618\ : Span12Mux_v
    port map (
            O => \N__42648\,
            I => \N__42637\
        );

    \I__9617\ : Span4Mux_h
    port map (
            O => \N__42643\,
            I => \N__42634\
        );

    \I__9616\ : LocalMux
    port map (
            O => \N__42640\,
            I => \N__42631\
        );

    \I__9615\ : Odrv12
    port map (
            O => \N__42637\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9614\ : Odrv4
    port map (
            O => \N__42634\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9613\ : Odrv4
    port map (
            O => \N__42631\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__9612\ : InMux
    port map (
            O => \N__42624\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__9611\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42617\
        );

    \I__9610\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42614\
        );

    \I__9609\ : LocalMux
    port map (
            O => \N__42617\,
            I => \N__42608\
        );

    \I__9608\ : LocalMux
    port map (
            O => \N__42614\,
            I => \N__42608\
        );

    \I__9607\ : InMux
    port map (
            O => \N__42613\,
            I => \N__42605\
        );

    \I__9606\ : Span4Mux_v
    port map (
            O => \N__42608\,
            I => \N__42599\
        );

    \I__9605\ : LocalMux
    port map (
            O => \N__42605\,
            I => \N__42599\
        );

    \I__9604\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42596\
        );

    \I__9603\ : Span4Mux_h
    port map (
            O => \N__42599\,
            I => \N__42593\
        );

    \I__9602\ : LocalMux
    port map (
            O => \N__42596\,
            I => \N__42590\
        );

    \I__9601\ : Odrv4
    port map (
            O => \N__42593\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9600\ : Odrv4
    port map (
            O => \N__42590\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__9599\ : InMux
    port map (
            O => \N__42585\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__9598\ : CascadeMux
    port map (
            O => \N__42582\,
            I => \N__42578\
        );

    \I__9597\ : InMux
    port map (
            O => \N__42581\,
            I => \N__42573\
        );

    \I__9596\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42568\
        );

    \I__9595\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42568\
        );

    \I__9594\ : InMux
    port map (
            O => \N__42576\,
            I => \N__42565\
        );

    \I__9593\ : LocalMux
    port map (
            O => \N__42573\,
            I => \N__42562\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__42568\,
            I => \N__42557\
        );

    \I__9591\ : LocalMux
    port map (
            O => \N__42565\,
            I => \N__42557\
        );

    \I__9590\ : Span4Mux_v
    port map (
            O => \N__42562\,
            I => \N__42554\
        );

    \I__9589\ : Span4Mux_v
    port map (
            O => \N__42557\,
            I => \N__42551\
        );

    \I__9588\ : Odrv4
    port map (
            O => \N__42554\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9587\ : Odrv4
    port map (
            O => \N__42551\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9586\ : InMux
    port map (
            O => \N__42546\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__9585\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42540\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__42540\,
            I => \N__42537\
        );

    \I__9583\ : Span4Mux_h
    port map (
            O => \N__42537\,
            I => \N__42534\
        );

    \I__9582\ : Odrv4
    port map (
            O => \N__42534\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__9581\ : InMux
    port map (
            O => \N__42531\,
            I => \N__42528\
        );

    \I__9580\ : LocalMux
    port map (
            O => \N__42528\,
            I => \N__42525\
        );

    \I__9579\ : Span4Mux_h
    port map (
            O => \N__42525\,
            I => \N__42522\
        );

    \I__9578\ : Odrv4
    port map (
            O => \N__42522\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__9577\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42516\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__42516\,
            I => \N__42513\
        );

    \I__9575\ : Span4Mux_h
    port map (
            O => \N__42513\,
            I => \N__42510\
        );

    \I__9574\ : Odrv4
    port map (
            O => \N__42510\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__9573\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42504\
        );

    \I__9572\ : LocalMux
    port map (
            O => \N__42504\,
            I => \N__42501\
        );

    \I__9571\ : Span4Mux_h
    port map (
            O => \N__42501\,
            I => \N__42498\
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__42498\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__9569\ : CascadeMux
    port map (
            O => \N__42495\,
            I => \N__42492\
        );

    \I__9568\ : InMux
    port map (
            O => \N__42492\,
            I => \N__42489\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__42489\,
            I => \N__42484\
        );

    \I__9566\ : InMux
    port map (
            O => \N__42488\,
            I => \N__42481\
        );

    \I__9565\ : InMux
    port map (
            O => \N__42487\,
            I => \N__42478\
        );

    \I__9564\ : Span4Mux_h
    port map (
            O => \N__42484\,
            I => \N__42473\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__42481\,
            I => \N__42473\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__42478\,
            I => \N__42469\
        );

    \I__9561\ : Span4Mux_h
    port map (
            O => \N__42473\,
            I => \N__42466\
        );

    \I__9560\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42463\
        );

    \I__9559\ : Odrv12
    port map (
            O => \N__42469\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9558\ : Odrv4
    port map (
            O => \N__42466\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__42463\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9556\ : InMux
    port map (
            O => \N__42456\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__9555\ : CascadeMux
    port map (
            O => \N__42453\,
            I => \N__42450\
        );

    \I__9554\ : InMux
    port map (
            O => \N__42450\,
            I => \N__42446\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42449\,
            I => \N__42442\
        );

    \I__9552\ : LocalMux
    port map (
            O => \N__42446\,
            I => \N__42439\
        );

    \I__9551\ : InMux
    port map (
            O => \N__42445\,
            I => \N__42436\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__42442\,
            I => \N__42431\
        );

    \I__9549\ : Span4Mux_h
    port map (
            O => \N__42439\,
            I => \N__42431\
        );

    \I__9548\ : LocalMux
    port map (
            O => \N__42436\,
            I => \N__42428\
        );

    \I__9547\ : Span4Mux_h
    port map (
            O => \N__42431\,
            I => \N__42424\
        );

    \I__9546\ : Span12Mux_h
    port map (
            O => \N__42428\,
            I => \N__42421\
        );

    \I__9545\ : InMux
    port map (
            O => \N__42427\,
            I => \N__42418\
        );

    \I__9544\ : Odrv4
    port map (
            O => \N__42424\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9543\ : Odrv12
    port map (
            O => \N__42421\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9542\ : LocalMux
    port map (
            O => \N__42418\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9541\ : InMux
    port map (
            O => \N__42411\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__9540\ : CascadeMux
    port map (
            O => \N__42408\,
            I => \N__42404\
        );

    \I__9539\ : InMux
    port map (
            O => \N__42407\,
            I => \N__42401\
        );

    \I__9538\ : InMux
    port map (
            O => \N__42404\,
            I => \N__42396\
        );

    \I__9537\ : LocalMux
    port map (
            O => \N__42401\,
            I => \N__42393\
        );

    \I__9536\ : InMux
    port map (
            O => \N__42400\,
            I => \N__42390\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42399\,
            I => \N__42387\
        );

    \I__9534\ : LocalMux
    port map (
            O => \N__42396\,
            I => \N__42382\
        );

    \I__9533\ : Span4Mux_h
    port map (
            O => \N__42393\,
            I => \N__42382\
        );

    \I__9532\ : LocalMux
    port map (
            O => \N__42390\,
            I => \N__42379\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__42387\,
            I => \N__42374\
        );

    \I__9530\ : Span4Mux_h
    port map (
            O => \N__42382\,
            I => \N__42374\
        );

    \I__9529\ : Span4Mux_v
    port map (
            O => \N__42379\,
            I => \N__42371\
        );

    \I__9528\ : Span4Mux_h
    port map (
            O => \N__42374\,
            I => \N__42368\
        );

    \I__9527\ : Odrv4
    port map (
            O => \N__42371\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__42368\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9525\ : InMux
    port map (
            O => \N__42363\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__9524\ : CascadeMux
    port map (
            O => \N__42360\,
            I => \N__42356\
        );

    \I__9523\ : CascadeMux
    port map (
            O => \N__42359\,
            I => \N__42353\
        );

    \I__9522\ : InMux
    port map (
            O => \N__42356\,
            I => \N__42350\
        );

    \I__9521\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42347\
        );

    \I__9520\ : LocalMux
    port map (
            O => \N__42350\,
            I => \N__42340\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__42347\,
            I => \N__42340\
        );

    \I__9518\ : InMux
    port map (
            O => \N__42346\,
            I => \N__42337\
        );

    \I__9517\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42334\
        );

    \I__9516\ : Span4Mux_v
    port map (
            O => \N__42340\,
            I => \N__42327\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__42337\,
            I => \N__42327\
        );

    \I__9514\ : LocalMux
    port map (
            O => \N__42334\,
            I => \N__42327\
        );

    \I__9513\ : Span4Mux_h
    port map (
            O => \N__42327\,
            I => \N__42324\
        );

    \I__9512\ : Odrv4
    port map (
            O => \N__42324\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42321\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__9510\ : CascadeMux
    port map (
            O => \N__42318\,
            I => \N__42315\
        );

    \I__9509\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42312\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42312\,
            I => \N__42309\
        );

    \I__9507\ : Span4Mux_h
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__9506\ : Odrv4
    port map (
            O => \N__42306\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__9505\ : InMux
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__42300\,
            I => \N__42297\
        );

    \I__9503\ : Span4Mux_h
    port map (
            O => \N__42297\,
            I => \N__42293\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42296\,
            I => \N__42290\
        );

    \I__9501\ : Odrv4
    port map (
            O => \N__42293\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42290\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__9499\ : InMux
    port map (
            O => \N__42285\,
            I => \N__42278\
        );

    \I__9498\ : InMux
    port map (
            O => \N__42284\,
            I => \N__42278\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42283\,
            I => \N__42274\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42278\,
            I => \N__42271\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42268\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__42274\,
            I => \N__42263\
        );

    \I__9493\ : Span4Mux_v
    port map (
            O => \N__42271\,
            I => \N__42263\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__42268\,
            I => \N__42260\
        );

    \I__9491\ : Odrv4
    port map (
            O => \N__42263\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9490\ : Odrv4
    port map (
            O => \N__42260\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__9489\ : CascadeMux
    port map (
            O => \N__42255\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42249\
        );

    \I__9487\ : LocalMux
    port map (
            O => \N__42249\,
            I => \N__42246\
        );

    \I__9486\ : Odrv4
    port map (
            O => \N__42246\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42243\,
            I => \N__42239\
        );

    \I__9484\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42236\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42239\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__9482\ : LocalMux
    port map (
            O => \N__42236\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__9481\ : InMux
    port map (
            O => \N__42231\,
            I => \N__42226\
        );

    \I__9480\ : InMux
    port map (
            O => \N__42230\,
            I => \N__42223\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42229\,
            I => \N__42220\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__42226\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42223\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9476\ : LocalMux
    port map (
            O => \N__42220\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9475\ : CascadeMux
    port map (
            O => \N__42213\,
            I => \N__42209\
        );

    \I__9474\ : CascadeMux
    port map (
            O => \N__42212\,
            I => \N__42206\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42209\,
            I => \N__42203\
        );

    \I__9472\ : InMux
    port map (
            O => \N__42206\,
            I => \N__42200\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42203\,
            I => \N__42195\
        );

    \I__9470\ : LocalMux
    port map (
            O => \N__42200\,
            I => \N__42195\
        );

    \I__9469\ : Odrv12
    port map (
            O => \N__42195\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__9468\ : InMux
    port map (
            O => \N__42192\,
            I => \N__42187\
        );

    \I__9467\ : InMux
    port map (
            O => \N__42191\,
            I => \N__42184\
        );

    \I__9466\ : InMux
    port map (
            O => \N__42190\,
            I => \N__42181\
        );

    \I__9465\ : LocalMux
    port map (
            O => \N__42187\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9464\ : LocalMux
    port map (
            O => \N__42184\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__42181\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42174\,
            I => \N__42171\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42171\,
            I => \N__42168\
        );

    \I__9460\ : Span4Mux_h
    port map (
            O => \N__42168\,
            I => \N__42165\
        );

    \I__9459\ : Odrv4
    port map (
            O => \N__42165\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42162\,
            I => \N__42159\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42159\,
            I => \N__42156\
        );

    \I__9456\ : Odrv12
    port map (
            O => \N__42156\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__9455\ : InMux
    port map (
            O => \N__42153\,
            I => \N__42150\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__42150\,
            I => \N__42147\
        );

    \I__9453\ : Odrv4
    port map (
            O => \N__42147\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__9452\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42141\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__42141\,
            I => \N__42138\
        );

    \I__9450\ : Odrv4
    port map (
            O => \N__42138\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42132\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__42129\
        );

    \I__9447\ : Span4Mux_v
    port map (
            O => \N__42129\,
            I => \N__42126\
        );

    \I__9446\ : Odrv4
    port map (
            O => \N__42126\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__9445\ : IoInMux
    port map (
            O => \N__42123\,
            I => \N__42089\
        );

    \I__9444\ : InMux
    port map (
            O => \N__42122\,
            I => \N__42086\
        );

    \I__9443\ : InMux
    port map (
            O => \N__42121\,
            I => \N__42079\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42120\,
            I => \N__42079\
        );

    \I__9441\ : InMux
    port map (
            O => \N__42119\,
            I => \N__42079\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42118\,
            I => \N__42070\
        );

    \I__9439\ : InMux
    port map (
            O => \N__42117\,
            I => \N__42070\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42116\,
            I => \N__42070\
        );

    \I__9437\ : InMux
    port map (
            O => \N__42115\,
            I => \N__42070\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42114\,
            I => \N__42061\
        );

    \I__9435\ : InMux
    port map (
            O => \N__42113\,
            I => \N__42061\
        );

    \I__9434\ : InMux
    port map (
            O => \N__42112\,
            I => \N__42061\
        );

    \I__9433\ : InMux
    port map (
            O => \N__42111\,
            I => \N__42061\
        );

    \I__9432\ : InMux
    port map (
            O => \N__42110\,
            I => \N__42052\
        );

    \I__9431\ : InMux
    port map (
            O => \N__42109\,
            I => \N__42052\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42108\,
            I => \N__42052\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42107\,
            I => \N__42052\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42106\,
            I => \N__42043\
        );

    \I__9427\ : InMux
    port map (
            O => \N__42105\,
            I => \N__42043\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42104\,
            I => \N__42043\
        );

    \I__9425\ : InMux
    port map (
            O => \N__42103\,
            I => \N__42043\
        );

    \I__9424\ : InMux
    port map (
            O => \N__42102\,
            I => \N__42034\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42101\,
            I => \N__42034\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42100\,
            I => \N__42034\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42034\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42098\,
            I => \N__42027\
        );

    \I__9419\ : InMux
    port map (
            O => \N__42097\,
            I => \N__42027\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42027\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42095\,
            I => \N__42018\
        );

    \I__9416\ : InMux
    port map (
            O => \N__42094\,
            I => \N__42018\
        );

    \I__9415\ : InMux
    port map (
            O => \N__42093\,
            I => \N__42018\
        );

    \I__9414\ : InMux
    port map (
            O => \N__42092\,
            I => \N__42018\
        );

    \I__9413\ : LocalMux
    port map (
            O => \N__42089\,
            I => \N__42015\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__42086\,
            I => \N__42012\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42079\,
            I => \N__42007\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__42070\,
            I => \N__42007\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__42061\,
            I => \N__42002\
        );

    \I__9408\ : LocalMux
    port map (
            O => \N__42052\,
            I => \N__42002\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42043\,
            I => \N__41997\
        );

    \I__9406\ : LocalMux
    port map (
            O => \N__42034\,
            I => \N__41997\
        );

    \I__9405\ : LocalMux
    port map (
            O => \N__42027\,
            I => \N__41992\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__42018\,
            I => \N__41992\
        );

    \I__9403\ : IoSpan4Mux
    port map (
            O => \N__42015\,
            I => \N__41989\
        );

    \I__9402\ : Span4Mux_h
    port map (
            O => \N__42012\,
            I => \N__41984\
        );

    \I__9401\ : Span4Mux_h
    port map (
            O => \N__42007\,
            I => \N__41984\
        );

    \I__9400\ : Span4Mux_h
    port map (
            O => \N__42002\,
            I => \N__41981\
        );

    \I__9399\ : Span4Mux_h
    port map (
            O => \N__41997\,
            I => \N__41978\
        );

    \I__9398\ : Span12Mux_s10_h
    port map (
            O => \N__41992\,
            I => \N__41975\
        );

    \I__9397\ : Span4Mux_s1_v
    port map (
            O => \N__41989\,
            I => \N__41970\
        );

    \I__9396\ : Span4Mux_v
    port map (
            O => \N__41984\,
            I => \N__41970\
        );

    \I__9395\ : Span4Mux_v
    port map (
            O => \N__41981\,
            I => \N__41967\
        );

    \I__9394\ : Odrv4
    port map (
            O => \N__41978\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9393\ : Odrv12
    port map (
            O => \N__41975\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__41970\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9391\ : Odrv4
    port map (
            O => \N__41967\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__9390\ : InMux
    port map (
            O => \N__41958\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__9389\ : InMux
    port map (
            O => \N__41955\,
            I => \N__41952\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__41952\,
            I => \N__41948\
        );

    \I__9387\ : CascadeMux
    port map (
            O => \N__41951\,
            I => \N__41945\
        );

    \I__9386\ : Span4Mux_h
    port map (
            O => \N__41948\,
            I => \N__41941\
        );

    \I__9385\ : InMux
    port map (
            O => \N__41945\,
            I => \N__41937\
        );

    \I__9384\ : InMux
    port map (
            O => \N__41944\,
            I => \N__41934\
        );

    \I__9383\ : Sp12to4
    port map (
            O => \N__41941\,
            I => \N__41931\
        );

    \I__9382\ : InMux
    port map (
            O => \N__41940\,
            I => \N__41928\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__41937\,
            I => \N__41924\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__41934\,
            I => \N__41921\
        );

    \I__9379\ : Span12Mux_v
    port map (
            O => \N__41931\,
            I => \N__41918\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41915\
        );

    \I__9377\ : InMux
    port map (
            O => \N__41927\,
            I => \N__41912\
        );

    \I__9376\ : Span4Mux_v
    port map (
            O => \N__41924\,
            I => \N__41909\
        );

    \I__9375\ : Span12Mux_v
    port map (
            O => \N__41921\,
            I => \N__41904\
        );

    \I__9374\ : Span12Mux_v
    port map (
            O => \N__41918\,
            I => \N__41904\
        );

    \I__9373\ : Span4Mux_h
    port map (
            O => \N__41915\,
            I => \N__41901\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__41912\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9371\ : Odrv4
    port map (
            O => \N__41909\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9370\ : Odrv12
    port map (
            O => \N__41904\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9369\ : Odrv4
    port map (
            O => \N__41901\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__9368\ : IoInMux
    port map (
            O => \N__41892\,
            I => \N__41889\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__41889\,
            I => \N__41886\
        );

    \I__9366\ : Span12Mux_s8_v
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__9365\ : Span12Mux_v
    port map (
            O => \N__41883\,
            I => \N__41879\
        );

    \I__9364\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41876\
        );

    \I__9363\ : Odrv12
    port map (
            O => \N__41879\,
            I => \T23_c\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__41876\,
            I => \T23_c\
        );

    \I__9361\ : InMux
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__41868\,
            I => \N__41864\
        );

    \I__9359\ : InMux
    port map (
            O => \N__41867\,
            I => \N__41861\
        );

    \I__9358\ : Span4Mux_v
    port map (
            O => \N__41864\,
            I => \N__41858\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__41861\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__9356\ : Odrv4
    port map (
            O => \N__41858\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__9355\ : CascadeMux
    port map (
            O => \N__41853\,
            I => \N__41850\
        );

    \I__9354\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41847\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__9352\ : Span4Mux_v
    port map (
            O => \N__41844\,
            I => \N__41841\
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__41841\,
            I => \phase_controller_inst2.stoper_tr.un4_running_df30\
        );

    \I__9350\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41835\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__41835\,
            I => \N__41829\
        );

    \I__9348\ : InMux
    port map (
            O => \N__41834\,
            I => \N__41824\
        );

    \I__9347\ : InMux
    port map (
            O => \N__41833\,
            I => \N__41824\
        );

    \I__9346\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41821\
        );

    \I__9345\ : Span4Mux_v
    port map (
            O => \N__41829\,
            I => \N__41818\
        );

    \I__9344\ : LocalMux
    port map (
            O => \N__41824\,
            I => \N__41815\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__41821\,
            I => \N__41812\
        );

    \I__9342\ : Odrv4
    port map (
            O => \N__41818\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9341\ : Odrv4
    port map (
            O => \N__41815\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9340\ : Odrv4
    port map (
            O => \N__41812\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__9339\ : InMux
    port map (
            O => \N__41805\,
            I => \N__41802\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__9337\ : Span4Mux_v
    port map (
            O => \N__41799\,
            I => \N__41795\
        );

    \I__9336\ : InMux
    port map (
            O => \N__41798\,
            I => \N__41792\
        );

    \I__9335\ : Odrv4
    port map (
            O => \N__41795\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__41792\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__9333\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41778\
        );

    \I__9332\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41778\
        );

    \I__9331\ : InMux
    port map (
            O => \N__41785\,
            I => \N__41778\
        );

    \I__9330\ : LocalMux
    port map (
            O => \N__41778\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__9329\ : InMux
    port map (
            O => \N__41775\,
            I => \N__41769\
        );

    \I__9328\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41762\
        );

    \I__9327\ : InMux
    port map (
            O => \N__41773\,
            I => \N__41762\
        );

    \I__9326\ : InMux
    port map (
            O => \N__41772\,
            I => \N__41762\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__41769\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__9324\ : LocalMux
    port map (
            O => \N__41762\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__9323\ : CascadeMux
    port map (
            O => \N__41757\,
            I => \N__41752\
        );

    \I__9322\ : CascadeMux
    port map (
            O => \N__41756\,
            I => \N__41749\
        );

    \I__9321\ : InMux
    port map (
            O => \N__41755\,
            I => \N__41745\
        );

    \I__9320\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41738\
        );

    \I__9319\ : InMux
    port map (
            O => \N__41749\,
            I => \N__41738\
        );

    \I__9318\ : InMux
    port map (
            O => \N__41748\,
            I => \N__41738\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__41745\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__41738\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__9315\ : CascadeMux
    port map (
            O => \N__41733\,
            I => \N__41730\
        );

    \I__9314\ : InMux
    port map (
            O => \N__41730\,
            I => \N__41727\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__41727\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__9312\ : CascadeMux
    port map (
            O => \N__41724\,
            I => \N__41720\
        );

    \I__9311\ : InMux
    port map (
            O => \N__41723\,
            I => \N__41712\
        );

    \I__9310\ : InMux
    port map (
            O => \N__41720\,
            I => \N__41712\
        );

    \I__9309\ : InMux
    port map (
            O => \N__41719\,
            I => \N__41712\
        );

    \I__9308\ : LocalMux
    port map (
            O => \N__41712\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__9307\ : InMux
    port map (
            O => \N__41709\,
            I => \N__41704\
        );

    \I__9306\ : InMux
    port map (
            O => \N__41708\,
            I => \N__41699\
        );

    \I__9305\ : InMux
    port map (
            O => \N__41707\,
            I => \N__41699\
        );

    \I__9304\ : LocalMux
    port map (
            O => \N__41704\,
            I => \N__41693\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__41699\,
            I => \N__41693\
        );

    \I__9302\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41690\
        );

    \I__9301\ : Span4Mux_h
    port map (
            O => \N__41693\,
            I => \N__41685\
        );

    \I__9300\ : LocalMux
    port map (
            O => \N__41690\,
            I => \N__41685\
        );

    \I__9299\ : Odrv4
    port map (
            O => \N__41685\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__9298\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41679\
        );

    \I__9297\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41675\
        );

    \I__9296\ : InMux
    port map (
            O => \N__41678\,
            I => \N__41672\
        );

    \I__9295\ : Odrv4
    port map (
            O => \N__41675\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__41672\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__9293\ : InMux
    port map (
            O => \N__41667\,
            I => \N__41664\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__41664\,
            I => \N__41661\
        );

    \I__9291\ : Odrv4
    port map (
            O => \N__41661\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__9290\ : InMux
    port map (
            O => \N__41658\,
            I => \N__41651\
        );

    \I__9289\ : InMux
    port map (
            O => \N__41657\,
            I => \N__41651\
        );

    \I__9288\ : InMux
    port map (
            O => \N__41656\,
            I => \N__41648\
        );

    \I__9287\ : LocalMux
    port map (
            O => \N__41651\,
            I => \N__41645\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__41648\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__9285\ : Odrv4
    port map (
            O => \N__41645\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__9284\ : InMux
    port map (
            O => \N__41640\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__9283\ : CascadeMux
    port map (
            O => \N__41637\,
            I => \N__41634\
        );

    \I__9282\ : InMux
    port map (
            O => \N__41634\,
            I => \N__41627\
        );

    \I__9281\ : InMux
    port map (
            O => \N__41633\,
            I => \N__41627\
        );

    \I__9280\ : InMux
    port map (
            O => \N__41632\,
            I => \N__41624\
        );

    \I__9279\ : LocalMux
    port map (
            O => \N__41627\,
            I => \N__41621\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__41624\,
            I => \N__41616\
        );

    \I__9277\ : Span4Mux_v
    port map (
            O => \N__41621\,
            I => \N__41616\
        );

    \I__9276\ : Odrv4
    port map (
            O => \N__41616\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__9275\ : InMux
    port map (
            O => \N__41613\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__9274\ : InMux
    port map (
            O => \N__41610\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__9273\ : InMux
    port map (
            O => \N__41607\,
            I => \bfn_17_10_0_\
        );

    \I__9272\ : InMux
    port map (
            O => \N__41604\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__9271\ : InMux
    port map (
            O => \N__41601\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__9270\ : InMux
    port map (
            O => \N__41598\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__9269\ : InMux
    port map (
            O => \N__41595\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__9268\ : InMux
    port map (
            O => \N__41592\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__9267\ : InMux
    port map (
            O => \N__41589\,
            I => \N__41585\
        );

    \I__9266\ : InMux
    port map (
            O => \N__41588\,
            I => \N__41582\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__41585\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__41582\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__9263\ : InMux
    port map (
            O => \N__41577\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__9262\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41570\
        );

    \I__9261\ : InMux
    port map (
            O => \N__41573\,
            I => \N__41567\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__41570\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__41567\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__9258\ : InMux
    port map (
            O => \N__41562\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__9257\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41555\
        );

    \I__9256\ : InMux
    port map (
            O => \N__41558\,
            I => \N__41552\
        );

    \I__9255\ : LocalMux
    port map (
            O => \N__41555\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__41552\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__9253\ : InMux
    port map (
            O => \N__41547\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__9252\ : InMux
    port map (
            O => \N__41544\,
            I => \N__41537\
        );

    \I__9251\ : InMux
    port map (
            O => \N__41543\,
            I => \N__41537\
        );

    \I__9250\ : InMux
    port map (
            O => \N__41542\,
            I => \N__41534\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__41537\,
            I => \N__41531\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__41534\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9247\ : Odrv4
    port map (
            O => \N__41531\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__9246\ : InMux
    port map (
            O => \N__41526\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__9245\ : CascadeMux
    port map (
            O => \N__41523\,
            I => \N__41519\
        );

    \I__9244\ : InMux
    port map (
            O => \N__41522\,
            I => \N__41514\
        );

    \I__9243\ : InMux
    port map (
            O => \N__41519\,
            I => \N__41514\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__41514\,
            I => \N__41510\
        );

    \I__9241\ : InMux
    port map (
            O => \N__41513\,
            I => \N__41507\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__41510\,
            I => \N__41504\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__41507\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9238\ : Odrv4
    port map (
            O => \N__41504\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__9237\ : InMux
    port map (
            O => \N__41499\,
            I => \bfn_17_9_0_\
        );

    \I__9236\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41489\
        );

    \I__9235\ : InMux
    port map (
            O => \N__41495\,
            I => \N__41489\
        );

    \I__9234\ : InMux
    port map (
            O => \N__41494\,
            I => \N__41486\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__41489\,
            I => \N__41483\
        );

    \I__9232\ : LocalMux
    port map (
            O => \N__41486\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__41483\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__9230\ : InMux
    port map (
            O => \N__41478\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__9229\ : CascadeMux
    port map (
            O => \N__41475\,
            I => \N__41472\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41472\,
            I => \N__41465\
        );

    \I__9227\ : InMux
    port map (
            O => \N__41471\,
            I => \N__41465\
        );

    \I__9226\ : InMux
    port map (
            O => \N__41470\,
            I => \N__41462\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__41465\,
            I => \N__41459\
        );

    \I__9224\ : LocalMux
    port map (
            O => \N__41462\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9223\ : Odrv4
    port map (
            O => \N__41459\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__9222\ : InMux
    port map (
            O => \N__41454\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__9221\ : InMux
    port map (
            O => \N__41451\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__9220\ : InMux
    port map (
            O => \N__41448\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__9219\ : InMux
    port map (
            O => \N__41445\,
            I => \N__41441\
        );

    \I__9218\ : InMux
    port map (
            O => \N__41444\,
            I => \N__41438\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__41441\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__41438\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41433\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__9214\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41427\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41423\
        );

    \I__9212\ : InMux
    port map (
            O => \N__41426\,
            I => \N__41420\
        );

    \I__9211\ : Span4Mux_v
    port map (
            O => \N__41423\,
            I => \N__41417\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41420\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9209\ : Odrv4
    port map (
            O => \N__41417\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41412\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41409\,
            I => \N__41405\
        );

    \I__9206\ : InMux
    port map (
            O => \N__41408\,
            I => \N__41402\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41405\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9204\ : LocalMux
    port map (
            O => \N__41402\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__9203\ : InMux
    port map (
            O => \N__41397\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41394\,
            I => \N__41390\
        );

    \I__9201\ : InMux
    port map (
            O => \N__41393\,
            I => \N__41387\
        );

    \I__9200\ : LocalMux
    port map (
            O => \N__41390\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__41387\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__9198\ : InMux
    port map (
            O => \N__41382\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41375\
        );

    \I__9196\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41372\
        );

    \I__9195\ : LocalMux
    port map (
            O => \N__41375\,
            I => \N__41369\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__41372\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9193\ : Odrv4
    port map (
            O => \N__41369\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__9192\ : InMux
    port map (
            O => \N__41364\,
            I => \bfn_17_8_0_\
        );

    \I__9191\ : InMux
    port map (
            O => \N__41361\,
            I => \N__41357\
        );

    \I__9190\ : InMux
    port map (
            O => \N__41360\,
            I => \N__41354\
        );

    \I__9189\ : LocalMux
    port map (
            O => \N__41357\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41354\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41349\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__9186\ : InMux
    port map (
            O => \N__41346\,
            I => \N__41342\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41345\,
            I => \N__41339\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__41342\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__41339\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__9182\ : InMux
    port map (
            O => \N__41334\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41331\,
            I => \N__41327\
        );

    \I__9180\ : InMux
    port map (
            O => \N__41330\,
            I => \N__41324\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__41327\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__41324\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__9177\ : InMux
    port map (
            O => \N__41319\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41316\,
            I => \N__41313\
        );

    \I__9175\ : LocalMux
    port map (
            O => \N__41313\,
            I => \N__41310\
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__41310\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9173\ : InMux
    port map (
            O => \N__41307\,
            I => \N__41303\
        );

    \I__9172\ : InMux
    port map (
            O => \N__41306\,
            I => \N__41298\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__41303\,
            I => \N__41295\
        );

    \I__9170\ : InMux
    port map (
            O => \N__41302\,
            I => \N__41290\
        );

    \I__9169\ : InMux
    port map (
            O => \N__41301\,
            I => \N__41290\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__41298\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9167\ : Odrv12
    port map (
            O => \N__41295\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__41290\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__9165\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41274\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41282\,
            I => \N__41274\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41281\,
            I => \N__41271\
        );

    \I__9162\ : InMux
    port map (
            O => \N__41280\,
            I => \N__41266\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41279\,
            I => \N__41266\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41274\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__41271\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__9158\ : LocalMux
    port map (
            O => \N__41266\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__9157\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41255\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41258\,
            I => \N__41252\
        );

    \I__9155\ : LocalMux
    port map (
            O => \N__41255\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41252\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41244\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__41244\,
            I => \N__41239\
        );

    \I__9151\ : InMux
    port map (
            O => \N__41243\,
            I => \N__41236\
        );

    \I__9150\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41232\
        );

    \I__9149\ : Span4Mux_v
    port map (
            O => \N__41239\,
            I => \N__41229\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41236\,
            I => \N__41226\
        );

    \I__9147\ : InMux
    port map (
            O => \N__41235\,
            I => \N__41223\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41232\,
            I => \N__41220\
        );

    \I__9145\ : Sp12to4
    port map (
            O => \N__41229\,
            I => \N__41217\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__41226\,
            I => \N__41212\
        );

    \I__9143\ : LocalMux
    port map (
            O => \N__41223\,
            I => \N__41212\
        );

    \I__9142\ : Span4Mux_h
    port map (
            O => \N__41220\,
            I => \N__41209\
        );

    \I__9141\ : Span12Mux_h
    port map (
            O => \N__41217\,
            I => \N__41206\
        );

    \I__9140\ : Span4Mux_h
    port map (
            O => \N__41212\,
            I => \N__41203\
        );

    \I__9139\ : Odrv4
    port map (
            O => \N__41209\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9138\ : Odrv12
    port map (
            O => \N__41206\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9137\ : Odrv4
    port map (
            O => \N__41203\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41193\
        );

    \I__9135\ : LocalMux
    port map (
            O => \N__41193\,
            I => \N__41156\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41192\,
            I => \N__41147\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41191\,
            I => \N__41147\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41190\,
            I => \N__41147\
        );

    \I__9131\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41147\
        );

    \I__9130\ : InMux
    port map (
            O => \N__41188\,
            I => \N__41144\
        );

    \I__9129\ : CascadeMux
    port map (
            O => \N__41187\,
            I => \N__41139\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41186\,
            I => \N__41129\
        );

    \I__9127\ : CascadeMux
    port map (
            O => \N__41185\,
            I => \N__41116\
        );

    \I__9126\ : InMux
    port map (
            O => \N__41184\,
            I => \N__41112\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41183\,
            I => \N__41106\
        );

    \I__9124\ : InMux
    port map (
            O => \N__41182\,
            I => \N__41099\
        );

    \I__9123\ : InMux
    port map (
            O => \N__41181\,
            I => \N__41099\
        );

    \I__9122\ : InMux
    port map (
            O => \N__41180\,
            I => \N__41087\
        );

    \I__9121\ : InMux
    port map (
            O => \N__41179\,
            I => \N__41087\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41178\,
            I => \N__41078\
        );

    \I__9119\ : InMux
    port map (
            O => \N__41177\,
            I => \N__41078\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41176\,
            I => \N__41078\
        );

    \I__9117\ : InMux
    port map (
            O => \N__41175\,
            I => \N__41078\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41174\,
            I => \N__41069\
        );

    \I__9115\ : InMux
    port map (
            O => \N__41173\,
            I => \N__41069\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41172\,
            I => \N__41069\
        );

    \I__9113\ : InMux
    port map (
            O => \N__41171\,
            I => \N__41069\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41066\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41063\
        );

    \I__9110\ : InMux
    port map (
            O => \N__41168\,
            I => \N__41060\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41167\,
            I => \N__41057\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41050\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41165\,
            I => \N__41050\
        );

    \I__9106\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41050\
        );

    \I__9105\ : InMux
    port map (
            O => \N__41163\,
            I => \N__41045\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41162\,
            I => \N__41045\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41161\,
            I => \N__41038\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41160\,
            I => \N__41038\
        );

    \I__9101\ : InMux
    port map (
            O => \N__41159\,
            I => \N__41038\
        );

    \I__9100\ : Span4Mux_h
    port map (
            O => \N__41156\,
            I => \N__41031\
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__41147\,
            I => \N__41031\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__41144\,
            I => \N__41031\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41143\,
            I => \N__41024\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41142\,
            I => \N__41024\
        );

    \I__9095\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41024\
        );

    \I__9094\ : InMux
    port map (
            O => \N__41138\,
            I => \N__41021\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41137\,
            I => \N__41018\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41136\,
            I => \N__41011\
        );

    \I__9091\ : InMux
    port map (
            O => \N__41135\,
            I => \N__41011\
        );

    \I__9090\ : InMux
    port map (
            O => \N__41134\,
            I => \N__41011\
        );

    \I__9089\ : InMux
    port map (
            O => \N__41133\,
            I => \N__41006\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41132\,
            I => \N__41006\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41129\,
            I => \N__41003\
        );

    \I__9086\ : InMux
    port map (
            O => \N__41128\,
            I => \N__40973\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41127\,
            I => \N__40973\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41126\,
            I => \N__40973\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41125\,
            I => \N__40973\
        );

    \I__9082\ : InMux
    port map (
            O => \N__41124\,
            I => \N__40973\
        );

    \I__9081\ : InMux
    port map (
            O => \N__41123\,
            I => \N__40973\
        );

    \I__9080\ : InMux
    port map (
            O => \N__41122\,
            I => \N__40973\
        );

    \I__9079\ : InMux
    port map (
            O => \N__41121\,
            I => \N__40973\
        );

    \I__9078\ : InMux
    port map (
            O => \N__41120\,
            I => \N__40964\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41119\,
            I => \N__40964\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41116\,
            I => \N__40964\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41115\,
            I => \N__40964\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41112\,
            I => \N__40961\
        );

    \I__9073\ : CascadeMux
    port map (
            O => \N__41111\,
            I => \N__40958\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41110\,
            I => \N__40941\
        );

    \I__9071\ : InMux
    port map (
            O => \N__41109\,
            I => \N__40941\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__40938\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41105\,
            I => \N__40933\
        );

    \I__9068\ : InMux
    port map (
            O => \N__41104\,
            I => \N__40933\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__41099\,
            I => \N__40930\
        );

    \I__9066\ : InMux
    port map (
            O => \N__41098\,
            I => \N__40919\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41097\,
            I => \N__40919\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41096\,
            I => \N__40919\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41095\,
            I => \N__40919\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41094\,
            I => \N__40919\
        );

    \I__9061\ : InMux
    port map (
            O => \N__41093\,
            I => \N__40914\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41092\,
            I => \N__40914\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__41087\,
            I => \N__40905\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41078\,
            I => \N__40905\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__41069\,
            I => \N__40905\
        );

    \I__9056\ : LocalMux
    port map (
            O => \N__41066\,
            I => \N__40905\
        );

    \I__9055\ : LocalMux
    port map (
            O => \N__41063\,
            I => \N__40902\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__41060\,
            I => \N__40899\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__41057\,
            I => \N__40886\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41050\,
            I => \N__40886\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__41045\,
            I => \N__40886\
        );

    \I__9050\ : LocalMux
    port map (
            O => \N__41038\,
            I => \N__40886\
        );

    \I__9049\ : Span4Mux_v
    port map (
            O => \N__41031\,
            I => \N__40886\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__41024\,
            I => \N__40886\
        );

    \I__9047\ : LocalMux
    port map (
            O => \N__41021\,
            I => \N__40881\
        );

    \I__9046\ : LocalMux
    port map (
            O => \N__41018\,
            I => \N__40881\
        );

    \I__9045\ : LocalMux
    port map (
            O => \N__41011\,
            I => \N__40876\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__41006\,
            I => \N__40876\
        );

    \I__9043\ : Span4Mux_v
    port map (
            O => \N__41003\,
            I => \N__40873\
        );

    \I__9042\ : InMux
    port map (
            O => \N__41002\,
            I => \N__40870\
        );

    \I__9041\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40857\
        );

    \I__9040\ : InMux
    port map (
            O => \N__41000\,
            I => \N__40857\
        );

    \I__9039\ : InMux
    port map (
            O => \N__40999\,
            I => \N__40857\
        );

    \I__9038\ : InMux
    port map (
            O => \N__40998\,
            I => \N__40857\
        );

    \I__9037\ : InMux
    port map (
            O => \N__40997\,
            I => \N__40857\
        );

    \I__9036\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40857\
        );

    \I__9035\ : InMux
    port map (
            O => \N__40995\,
            I => \N__40844\
        );

    \I__9034\ : InMux
    port map (
            O => \N__40994\,
            I => \N__40844\
        );

    \I__9033\ : InMux
    port map (
            O => \N__40993\,
            I => \N__40844\
        );

    \I__9032\ : InMux
    port map (
            O => \N__40992\,
            I => \N__40844\
        );

    \I__9031\ : InMux
    port map (
            O => \N__40991\,
            I => \N__40844\
        );

    \I__9030\ : InMux
    port map (
            O => \N__40990\,
            I => \N__40844\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__40973\,
            I => \N__40837\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__40964\,
            I => \N__40837\
        );

    \I__9027\ : Span4Mux_h
    port map (
            O => \N__40961\,
            I => \N__40837\
        );

    \I__9026\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40828\
        );

    \I__9025\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40828\
        );

    \I__9024\ : InMux
    port map (
            O => \N__40956\,
            I => \N__40828\
        );

    \I__9023\ : InMux
    port map (
            O => \N__40955\,
            I => \N__40828\
        );

    \I__9022\ : InMux
    port map (
            O => \N__40954\,
            I => \N__40821\
        );

    \I__9021\ : InMux
    port map (
            O => \N__40953\,
            I => \N__40821\
        );

    \I__9020\ : InMux
    port map (
            O => \N__40952\,
            I => \N__40821\
        );

    \I__9019\ : InMux
    port map (
            O => \N__40951\,
            I => \N__40814\
        );

    \I__9018\ : InMux
    port map (
            O => \N__40950\,
            I => \N__40814\
        );

    \I__9017\ : InMux
    port map (
            O => \N__40949\,
            I => \N__40814\
        );

    \I__9016\ : InMux
    port map (
            O => \N__40948\,
            I => \N__40807\
        );

    \I__9015\ : InMux
    port map (
            O => \N__40947\,
            I => \N__40807\
        );

    \I__9014\ : InMux
    port map (
            O => \N__40946\,
            I => \N__40807\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__40941\,
            I => \N__40798\
        );

    \I__9012\ : Span4Mux_v
    port map (
            O => \N__40938\,
            I => \N__40798\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__40933\,
            I => \N__40798\
        );

    \I__9010\ : Span4Mux_h
    port map (
            O => \N__40930\,
            I => \N__40798\
        );

    \I__9009\ : LocalMux
    port map (
            O => \N__40919\,
            I => \N__40789\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__40914\,
            I => \N__40789\
        );

    \I__9007\ : Sp12to4
    port map (
            O => \N__40905\,
            I => \N__40789\
        );

    \I__9006\ : Span12Mux_s10_h
    port map (
            O => \N__40902\,
            I => \N__40789\
        );

    \I__9005\ : Span4Mux_v
    port map (
            O => \N__40899\,
            I => \N__40778\
        );

    \I__9004\ : Span4Mux_v
    port map (
            O => \N__40886\,
            I => \N__40778\
        );

    \I__9003\ : Span4Mux_v
    port map (
            O => \N__40881\,
            I => \N__40778\
        );

    \I__9002\ : Span4Mux_h
    port map (
            O => \N__40876\,
            I => \N__40778\
        );

    \I__9001\ : Span4Mux_h
    port map (
            O => \N__40873\,
            I => \N__40778\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__40870\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__40857\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__40844\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8997\ : Odrv4
    port map (
            O => \N__40837\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__40828\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__40821\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8994\ : LocalMux
    port map (
            O => \N__40814\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__40807\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8992\ : Odrv4
    port map (
            O => \N__40798\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8991\ : Odrv12
    port map (
            O => \N__40789\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8990\ : Odrv4
    port map (
            O => \N__40778\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__8989\ : InMux
    port map (
            O => \N__40755\,
            I => \N__40752\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__40752\,
            I => \N__40748\
        );

    \I__8987\ : InMux
    port map (
            O => \N__40751\,
            I => \N__40745\
        );

    \I__8986\ : Span4Mux_h
    port map (
            O => \N__40748\,
            I => \N__40742\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__40745\,
            I => \N__40739\
        );

    \I__8984\ : Span4Mux_h
    port map (
            O => \N__40742\,
            I => \N__40735\
        );

    \I__8983\ : Span4Mux_h
    port map (
            O => \N__40739\,
            I => \N__40732\
        );

    \I__8982\ : InMux
    port map (
            O => \N__40738\,
            I => \N__40729\
        );

    \I__8981\ : Span4Mux_v
    port map (
            O => \N__40735\,
            I => \N__40726\
        );

    \I__8980\ : Span4Mux_h
    port map (
            O => \N__40732\,
            I => \N__40723\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__40729\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__40726\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__8977\ : Odrv4
    port map (
            O => \N__40723\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__8976\ : CascadeMux
    port map (
            O => \N__40716\,
            I => \N__40712\
        );

    \I__8975\ : InMux
    port map (
            O => \N__40715\,
            I => \N__40708\
        );

    \I__8974\ : InMux
    port map (
            O => \N__40712\,
            I => \N__40705\
        );

    \I__8973\ : InMux
    port map (
            O => \N__40711\,
            I => \N__40702\
        );

    \I__8972\ : LocalMux
    port map (
            O => \N__40708\,
            I => \N__40699\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__40705\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8970\ : LocalMux
    port map (
            O => \N__40702\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8969\ : Odrv4
    port map (
            O => \N__40699\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__40692\,
            I => \N__40689\
        );

    \I__8967\ : InMux
    port map (
            O => \N__40689\,
            I => \N__40686\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__40686\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__8965\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40679\
        );

    \I__8964\ : InMux
    port map (
            O => \N__40682\,
            I => \N__40676\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__40679\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__40676\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8961\ : InMux
    port map (
            O => \N__40671\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__8960\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40665\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__40665\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\
        );

    \I__8958\ : CascadeMux
    port map (
            O => \N__40662\,
            I => \N__40659\
        );

    \I__8957\ : InMux
    port map (
            O => \N__40659\,
            I => \N__40655\
        );

    \I__8956\ : InMux
    port map (
            O => \N__40658\,
            I => \N__40652\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__40655\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__40652\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8953\ : InMux
    port map (
            O => \N__40647\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__8952\ : InMux
    port map (
            O => \N__40644\,
            I => \N__40640\
        );

    \I__8951\ : InMux
    port map (
            O => \N__40643\,
            I => \N__40637\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__40640\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__40637\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8948\ : InMux
    port map (
            O => \N__40632\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__8947\ : InMux
    port map (
            O => \N__40629\,
            I => \N__40622\
        );

    \I__8946\ : CascadeMux
    port map (
            O => \N__40628\,
            I => \N__40618\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__40627\,
            I => \N__40591\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__40626\,
            I => \N__40588\
        );

    \I__8943\ : InMux
    port map (
            O => \N__40625\,
            I => \N__40567\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__40622\,
            I => \N__40561\
        );

    \I__8941\ : InMux
    port map (
            O => \N__40621\,
            I => \N__40544\
        );

    \I__8940\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40544\
        );

    \I__8939\ : InMux
    port map (
            O => \N__40617\,
            I => \N__40544\
        );

    \I__8938\ : InMux
    port map (
            O => \N__40616\,
            I => \N__40544\
        );

    \I__8937\ : InMux
    port map (
            O => \N__40615\,
            I => \N__40544\
        );

    \I__8936\ : InMux
    port map (
            O => \N__40614\,
            I => \N__40544\
        );

    \I__8935\ : InMux
    port map (
            O => \N__40613\,
            I => \N__40544\
        );

    \I__8934\ : InMux
    port map (
            O => \N__40612\,
            I => \N__40544\
        );

    \I__8933\ : InMux
    port map (
            O => \N__40611\,
            I => \N__40531\
        );

    \I__8932\ : InMux
    port map (
            O => \N__40610\,
            I => \N__40531\
        );

    \I__8931\ : InMux
    port map (
            O => \N__40609\,
            I => \N__40531\
        );

    \I__8930\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40531\
        );

    \I__8929\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40531\
        );

    \I__8928\ : InMux
    port map (
            O => \N__40606\,
            I => \N__40531\
        );

    \I__8927\ : InMux
    port map (
            O => \N__40605\,
            I => \N__40528\
        );

    \I__8926\ : InMux
    port map (
            O => \N__40604\,
            I => \N__40519\
        );

    \I__8925\ : InMux
    port map (
            O => \N__40603\,
            I => \N__40519\
        );

    \I__8924\ : InMux
    port map (
            O => \N__40602\,
            I => \N__40519\
        );

    \I__8923\ : InMux
    port map (
            O => \N__40601\,
            I => \N__40519\
        );

    \I__8922\ : InMux
    port map (
            O => \N__40600\,
            I => \N__40512\
        );

    \I__8921\ : InMux
    port map (
            O => \N__40599\,
            I => \N__40512\
        );

    \I__8920\ : InMux
    port map (
            O => \N__40598\,
            I => \N__40512\
        );

    \I__8919\ : InMux
    port map (
            O => \N__40597\,
            I => \N__40507\
        );

    \I__8918\ : InMux
    port map (
            O => \N__40596\,
            I => \N__40507\
        );

    \I__8917\ : InMux
    port map (
            O => \N__40595\,
            I => \N__40502\
        );

    \I__8916\ : InMux
    port map (
            O => \N__40594\,
            I => \N__40502\
        );

    \I__8915\ : InMux
    port map (
            O => \N__40591\,
            I => \N__40487\
        );

    \I__8914\ : InMux
    port map (
            O => \N__40588\,
            I => \N__40487\
        );

    \I__8913\ : InMux
    port map (
            O => \N__40587\,
            I => \N__40487\
        );

    \I__8912\ : InMux
    port map (
            O => \N__40586\,
            I => \N__40487\
        );

    \I__8911\ : InMux
    port map (
            O => \N__40585\,
            I => \N__40487\
        );

    \I__8910\ : InMux
    port map (
            O => \N__40584\,
            I => \N__40487\
        );

    \I__8909\ : InMux
    port map (
            O => \N__40583\,
            I => \N__40487\
        );

    \I__8908\ : InMux
    port map (
            O => \N__40582\,
            I => \N__40479\
        );

    \I__8907\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40476\
        );

    \I__8906\ : InMux
    port map (
            O => \N__40580\,
            I => \N__40473\
        );

    \I__8905\ : InMux
    port map (
            O => \N__40579\,
            I => \N__40466\
        );

    \I__8904\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40466\
        );

    \I__8903\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40466\
        );

    \I__8902\ : InMux
    port map (
            O => \N__40576\,
            I => \N__40453\
        );

    \I__8901\ : InMux
    port map (
            O => \N__40575\,
            I => \N__40453\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40574\,
            I => \N__40453\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40573\,
            I => \N__40453\
        );

    \I__8898\ : InMux
    port map (
            O => \N__40572\,
            I => \N__40453\
        );

    \I__8897\ : InMux
    port map (
            O => \N__40571\,
            I => \N__40453\
        );

    \I__8896\ : InMux
    port map (
            O => \N__40570\,
            I => \N__40438\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__40567\,
            I => \N__40435\
        );

    \I__8894\ : InMux
    port map (
            O => \N__40566\,
            I => \N__40428\
        );

    \I__8893\ : InMux
    port map (
            O => \N__40565\,
            I => \N__40428\
        );

    \I__8892\ : InMux
    port map (
            O => \N__40564\,
            I => \N__40428\
        );

    \I__8891\ : Span4Mux_h
    port map (
            O => \N__40561\,
            I => \N__40423\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__40544\,
            I => \N__40423\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__40531\,
            I => \N__40420\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__40528\,
            I => \N__40417\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__40519\,
            I => \N__40412\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__40512\,
            I => \N__40412\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__40507\,
            I => \N__40407\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__40502\,
            I => \N__40407\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__40487\,
            I => \N__40404\
        );

    \I__8882\ : InMux
    port map (
            O => \N__40486\,
            I => \N__40393\
        );

    \I__8881\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40393\
        );

    \I__8880\ : InMux
    port map (
            O => \N__40484\,
            I => \N__40393\
        );

    \I__8879\ : InMux
    port map (
            O => \N__40483\,
            I => \N__40393\
        );

    \I__8878\ : InMux
    port map (
            O => \N__40482\,
            I => \N__40393\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__40479\,
            I => \N__40388\
        );

    \I__8876\ : LocalMux
    port map (
            O => \N__40476\,
            I => \N__40388\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__40473\,
            I => \N__40381\
        );

    \I__8874\ : LocalMux
    port map (
            O => \N__40466\,
            I => \N__40381\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40453\,
            I => \N__40381\
        );

    \I__8872\ : InMux
    port map (
            O => \N__40452\,
            I => \N__40364\
        );

    \I__8871\ : InMux
    port map (
            O => \N__40451\,
            I => \N__40364\
        );

    \I__8870\ : InMux
    port map (
            O => \N__40450\,
            I => \N__40364\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40449\,
            I => \N__40364\
        );

    \I__8868\ : InMux
    port map (
            O => \N__40448\,
            I => \N__40364\
        );

    \I__8867\ : InMux
    port map (
            O => \N__40447\,
            I => \N__40364\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40446\,
            I => \N__40364\
        );

    \I__8865\ : InMux
    port map (
            O => \N__40445\,
            I => \N__40364\
        );

    \I__8864\ : InMux
    port map (
            O => \N__40444\,
            I => \N__40358\
        );

    \I__8863\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40351\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40442\,
            I => \N__40351\
        );

    \I__8861\ : InMux
    port map (
            O => \N__40441\,
            I => \N__40351\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__40438\,
            I => \N__40344\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__40435\,
            I => \N__40344\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__40428\,
            I => \N__40344\
        );

    \I__8857\ : Span4Mux_v
    port map (
            O => \N__40423\,
            I => \N__40339\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__40420\,
            I => \N__40339\
        );

    \I__8855\ : Span4Mux_v
    port map (
            O => \N__40417\,
            I => \N__40336\
        );

    \I__8854\ : Span4Mux_v
    port map (
            O => \N__40412\,
            I => \N__40333\
        );

    \I__8853\ : Span4Mux_h
    port map (
            O => \N__40407\,
            I => \N__40326\
        );

    \I__8852\ : Span4Mux_h
    port map (
            O => \N__40404\,
            I => \N__40326\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40393\,
            I => \N__40326\
        );

    \I__8850\ : Span4Mux_h
    port map (
            O => \N__40388\,
            I => \N__40319\
        );

    \I__8849\ : Span4Mux_v
    port map (
            O => \N__40381\,
            I => \N__40319\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__40364\,
            I => \N__40319\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40363\,
            I => \N__40312\
        );

    \I__8846\ : InMux
    port map (
            O => \N__40362\,
            I => \N__40312\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40361\,
            I => \N__40312\
        );

    \I__8844\ : LocalMux
    port map (
            O => \N__40358\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__40351\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8842\ : Odrv4
    port map (
            O => \N__40344\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8841\ : Odrv4
    port map (
            O => \N__40339\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8840\ : Odrv4
    port map (
            O => \N__40336\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8839\ : Odrv4
    port map (
            O => \N__40333\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__40326\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8837\ : Odrv4
    port map (
            O => \N__40319\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40312\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40293\,
            I => \N__40288\
        );

    \I__8834\ : InMux
    port map (
            O => \N__40292\,
            I => \N__40285\
        );

    \I__8833\ : InMux
    port map (
            O => \N__40291\,
            I => \N__40282\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__40288\,
            I => \N__40279\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__40285\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8830\ : LocalMux
    port map (
            O => \N__40282\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8829\ : Odrv12
    port map (
            O => \N__40279\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__8828\ : CascadeMux
    port map (
            O => \N__40272\,
            I => \N__40257\
        );

    \I__8827\ : CascadeMux
    port map (
            O => \N__40271\,
            I => \N__40253\
        );

    \I__8826\ : CascadeMux
    port map (
            O => \N__40270\,
            I => \N__40250\
        );

    \I__8825\ : CascadeMux
    port map (
            O => \N__40269\,
            I => \N__40247\
        );

    \I__8824\ : CascadeMux
    port map (
            O => \N__40268\,
            I => \N__40242\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__40267\,
            I => \N__40239\
        );

    \I__8822\ : CascadeMux
    port map (
            O => \N__40266\,
            I => \N__40225\
        );

    \I__8821\ : InMux
    port map (
            O => \N__40265\,
            I => \N__40218\
        );

    \I__8820\ : InMux
    port map (
            O => \N__40264\,
            I => \N__40218\
        );

    \I__8819\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40218\
        );

    \I__8818\ : InMux
    port map (
            O => \N__40262\,
            I => \N__40209\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40261\,
            I => \N__40209\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40260\,
            I => \N__40209\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40209\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__40256\,
            I => \N__40205\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40253\,
            I => \N__40192\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40250\,
            I => \N__40187\
        );

    \I__8811\ : InMux
    port map (
            O => \N__40247\,
            I => \N__40187\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40246\,
            I => \N__40182\
        );

    \I__8809\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40182\
        );

    \I__8808\ : InMux
    port map (
            O => \N__40242\,
            I => \N__40179\
        );

    \I__8807\ : InMux
    port map (
            O => \N__40239\,
            I => \N__40176\
        );

    \I__8806\ : CascadeMux
    port map (
            O => \N__40238\,
            I => \N__40171\
        );

    \I__8805\ : CascadeMux
    port map (
            O => \N__40237\,
            I => \N__40167\
        );

    \I__8804\ : CascadeMux
    port map (
            O => \N__40236\,
            I => \N__40164\
        );

    \I__8803\ : CascadeMux
    port map (
            O => \N__40235\,
            I => \N__40160\
        );

    \I__8802\ : CascadeMux
    port map (
            O => \N__40234\,
            I => \N__40157\
        );

    \I__8801\ : CascadeMux
    port map (
            O => \N__40233\,
            I => \N__40154\
        );

    \I__8800\ : CascadeMux
    port map (
            O => \N__40232\,
            I => \N__40151\
        );

    \I__8799\ : CascadeMux
    port map (
            O => \N__40231\,
            I => \N__40147\
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__40230\,
            I => \N__40130\
        );

    \I__8797\ : CascadeMux
    port map (
            O => \N__40229\,
            I => \N__40122\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40228\,
            I => \N__40115\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40225\,
            I => \N__40115\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40218\,
            I => \N__40106\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40209\,
            I => \N__40106\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40208\,
            I => \N__40101\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40205\,
            I => \N__40101\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40204\,
            I => \N__40086\
        );

    \I__8789\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40086\
        );

    \I__8788\ : InMux
    port map (
            O => \N__40202\,
            I => \N__40086\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40201\,
            I => \N__40086\
        );

    \I__8786\ : InMux
    port map (
            O => \N__40200\,
            I => \N__40086\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40199\,
            I => \N__40086\
        );

    \I__8784\ : InMux
    port map (
            O => \N__40198\,
            I => \N__40086\
        );

    \I__8783\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40079\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40196\,
            I => \N__40079\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40195\,
            I => \N__40079\
        );

    \I__8780\ : LocalMux
    port map (
            O => \N__40192\,
            I => \N__40076\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40187\,
            I => \N__40073\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40182\,
            I => \N__40066\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__40179\,
            I => \N__40066\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__40176\,
            I => \N__40066\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40175\,
            I => \N__40061\
        );

    \I__8774\ : InMux
    port map (
            O => \N__40174\,
            I => \N__40061\
        );

    \I__8773\ : InMux
    port map (
            O => \N__40171\,
            I => \N__40052\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40170\,
            I => \N__40052\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40167\,
            I => \N__40052\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40052\
        );

    \I__8769\ : InMux
    port map (
            O => \N__40163\,
            I => \N__40043\
        );

    \I__8768\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40043\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40157\,
            I => \N__40043\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40154\,
            I => \N__40043\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40151\,
            I => \N__40040\
        );

    \I__8764\ : InMux
    port map (
            O => \N__40150\,
            I => \N__40035\
        );

    \I__8763\ : InMux
    port map (
            O => \N__40147\,
            I => \N__40035\
        );

    \I__8762\ : CascadeMux
    port map (
            O => \N__40146\,
            I => \N__40030\
        );

    \I__8761\ : CascadeMux
    port map (
            O => \N__40145\,
            I => \N__40026\
        );

    \I__8760\ : CascadeMux
    port map (
            O => \N__40144\,
            I => \N__40022\
        );

    \I__8759\ : CascadeMux
    port map (
            O => \N__40143\,
            I => \N__40017\
        );

    \I__8758\ : CascadeMux
    port map (
            O => \N__40142\,
            I => \N__40013\
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__40141\,
            I => \N__40009\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__40140\,
            I => \N__40004\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__40139\,
            I => \N__40000\
        );

    \I__8754\ : CascadeMux
    port map (
            O => \N__40138\,
            I => \N__39996\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__40137\,
            I => \N__39992\
        );

    \I__8752\ : CascadeMux
    port map (
            O => \N__40136\,
            I => \N__39989\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__40135\,
            I => \N__39985\
        );

    \I__8750\ : CascadeMux
    port map (
            O => \N__40134\,
            I => \N__39981\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__40133\,
            I => \N__39977\
        );

    \I__8748\ : InMux
    port map (
            O => \N__40130\,
            I => \N__39962\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__40129\,
            I => \N__39959\
        );

    \I__8746\ : InMux
    port map (
            O => \N__40128\,
            I => \N__39939\
        );

    \I__8745\ : InMux
    port map (
            O => \N__40127\,
            I => \N__39939\
        );

    \I__8744\ : InMux
    port map (
            O => \N__40126\,
            I => \N__39939\
        );

    \I__8743\ : InMux
    port map (
            O => \N__40125\,
            I => \N__39939\
        );

    \I__8742\ : InMux
    port map (
            O => \N__40122\,
            I => \N__39939\
        );

    \I__8741\ : InMux
    port map (
            O => \N__40121\,
            I => \N__39939\
        );

    \I__8740\ : InMux
    port map (
            O => \N__40120\,
            I => \N__39939\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__40115\,
            I => \N__39936\
        );

    \I__8738\ : InMux
    port map (
            O => \N__40114\,
            I => \N__39927\
        );

    \I__8737\ : InMux
    port map (
            O => \N__40113\,
            I => \N__39927\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40112\,
            I => \N__39927\
        );

    \I__8735\ : InMux
    port map (
            O => \N__40111\,
            I => \N__39927\
        );

    \I__8734\ : Span4Mux_v
    port map (
            O => \N__40106\,
            I => \N__39918\
        );

    \I__8733\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__39918\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__40086\,
            I => \N__39918\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__40079\,
            I => \N__39918\
        );

    \I__8730\ : Span4Mux_v
    port map (
            O => \N__40076\,
            I => \N__39901\
        );

    \I__8729\ : Span4Mux_h
    port map (
            O => \N__40073\,
            I => \N__39901\
        );

    \I__8728\ : Span4Mux_v
    port map (
            O => \N__40066\,
            I => \N__39901\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__40061\,
            I => \N__39901\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40052\,
            I => \N__39901\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40043\,
            I => \N__39901\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__40040\,
            I => \N__39901\
        );

    \I__8723\ : LocalMux
    port map (
            O => \N__40035\,
            I => \N__39901\
        );

    \I__8722\ : InMux
    port map (
            O => \N__40034\,
            I => \N__39884\
        );

    \I__8721\ : InMux
    port map (
            O => \N__40033\,
            I => \N__39884\
        );

    \I__8720\ : InMux
    port map (
            O => \N__40030\,
            I => \N__39884\
        );

    \I__8719\ : InMux
    port map (
            O => \N__40029\,
            I => \N__39884\
        );

    \I__8718\ : InMux
    port map (
            O => \N__40026\,
            I => \N__39884\
        );

    \I__8717\ : InMux
    port map (
            O => \N__40025\,
            I => \N__39884\
        );

    \I__8716\ : InMux
    port map (
            O => \N__40022\,
            I => \N__39884\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40021\,
            I => \N__39884\
        );

    \I__8714\ : InMux
    port map (
            O => \N__40020\,
            I => \N__39869\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40017\,
            I => \N__39869\
        );

    \I__8712\ : InMux
    port map (
            O => \N__40016\,
            I => \N__39869\
        );

    \I__8711\ : InMux
    port map (
            O => \N__40013\,
            I => \N__39869\
        );

    \I__8710\ : InMux
    port map (
            O => \N__40012\,
            I => \N__39869\
        );

    \I__8709\ : InMux
    port map (
            O => \N__40009\,
            I => \N__39869\
        );

    \I__8708\ : InMux
    port map (
            O => \N__40008\,
            I => \N__39869\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40007\,
            I => \N__39852\
        );

    \I__8706\ : InMux
    port map (
            O => \N__40004\,
            I => \N__39852\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40003\,
            I => \N__39852\
        );

    \I__8704\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39852\
        );

    \I__8703\ : InMux
    port map (
            O => \N__39999\,
            I => \N__39852\
        );

    \I__8702\ : InMux
    port map (
            O => \N__39996\,
            I => \N__39852\
        );

    \I__8701\ : InMux
    port map (
            O => \N__39995\,
            I => \N__39852\
        );

    \I__8700\ : InMux
    port map (
            O => \N__39992\,
            I => \N__39852\
        );

    \I__8699\ : InMux
    port map (
            O => \N__39989\,
            I => \N__39835\
        );

    \I__8698\ : InMux
    port map (
            O => \N__39988\,
            I => \N__39835\
        );

    \I__8697\ : InMux
    port map (
            O => \N__39985\,
            I => \N__39835\
        );

    \I__8696\ : InMux
    port map (
            O => \N__39984\,
            I => \N__39835\
        );

    \I__8695\ : InMux
    port map (
            O => \N__39981\,
            I => \N__39835\
        );

    \I__8694\ : InMux
    port map (
            O => \N__39980\,
            I => \N__39835\
        );

    \I__8693\ : InMux
    port map (
            O => \N__39977\,
            I => \N__39835\
        );

    \I__8692\ : InMux
    port map (
            O => \N__39976\,
            I => \N__39835\
        );

    \I__8691\ : CascadeMux
    port map (
            O => \N__39975\,
            I => \N__39832\
        );

    \I__8690\ : CascadeMux
    port map (
            O => \N__39974\,
            I => \N__39828\
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__39973\,
            I => \N__39824\
        );

    \I__8688\ : CascadeMux
    port map (
            O => \N__39972\,
            I => \N__39820\
        );

    \I__8687\ : CascadeMux
    port map (
            O => \N__39971\,
            I => \N__39816\
        );

    \I__8686\ : CascadeMux
    port map (
            O => \N__39970\,
            I => \N__39812\
        );

    \I__8685\ : CascadeMux
    port map (
            O => \N__39969\,
            I => \N__39808\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__39968\,
            I => \N__39804\
        );

    \I__8683\ : CascadeMux
    port map (
            O => \N__39967\,
            I => \N__39796\
        );

    \I__8682\ : CascadeMux
    port map (
            O => \N__39966\,
            I => \N__39792\
        );

    \I__8681\ : CascadeMux
    port map (
            O => \N__39965\,
            I => \N__39788\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__39962\,
            I => \N__39782\
        );

    \I__8679\ : InMux
    port map (
            O => \N__39959\,
            I => \N__39779\
        );

    \I__8678\ : InMux
    port map (
            O => \N__39958\,
            I => \N__39768\
        );

    \I__8677\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39768\
        );

    \I__8676\ : InMux
    port map (
            O => \N__39956\,
            I => \N__39768\
        );

    \I__8675\ : InMux
    port map (
            O => \N__39955\,
            I => \N__39768\
        );

    \I__8674\ : InMux
    port map (
            O => \N__39954\,
            I => \N__39768\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__39939\,
            I => \N__39765\
        );

    \I__8672\ : Span4Mux_h
    port map (
            O => \N__39936\,
            I => \N__39758\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__39927\,
            I => \N__39758\
        );

    \I__8670\ : Span4Mux_v
    port map (
            O => \N__39918\,
            I => \N__39758\
        );

    \I__8669\ : Span4Mux_h
    port map (
            O => \N__39901\,
            I => \N__39747\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__39884\,
            I => \N__39747\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__39869\,
            I => \N__39747\
        );

    \I__8666\ : LocalMux
    port map (
            O => \N__39852\,
            I => \N__39747\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__39835\,
            I => \N__39747\
        );

    \I__8664\ : InMux
    port map (
            O => \N__39832\,
            I => \N__39730\
        );

    \I__8663\ : InMux
    port map (
            O => \N__39831\,
            I => \N__39730\
        );

    \I__8662\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39730\
        );

    \I__8661\ : InMux
    port map (
            O => \N__39827\,
            I => \N__39730\
        );

    \I__8660\ : InMux
    port map (
            O => \N__39824\,
            I => \N__39730\
        );

    \I__8659\ : InMux
    port map (
            O => \N__39823\,
            I => \N__39730\
        );

    \I__8658\ : InMux
    port map (
            O => \N__39820\,
            I => \N__39730\
        );

    \I__8657\ : InMux
    port map (
            O => \N__39819\,
            I => \N__39730\
        );

    \I__8656\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39713\
        );

    \I__8655\ : InMux
    port map (
            O => \N__39815\,
            I => \N__39713\
        );

    \I__8654\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39713\
        );

    \I__8653\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39713\
        );

    \I__8652\ : InMux
    port map (
            O => \N__39808\,
            I => \N__39713\
        );

    \I__8651\ : InMux
    port map (
            O => \N__39807\,
            I => \N__39713\
        );

    \I__8650\ : InMux
    port map (
            O => \N__39804\,
            I => \N__39713\
        );

    \I__8649\ : InMux
    port map (
            O => \N__39803\,
            I => \N__39713\
        );

    \I__8648\ : InMux
    port map (
            O => \N__39802\,
            I => \N__39706\
        );

    \I__8647\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39706\
        );

    \I__8646\ : InMux
    port map (
            O => \N__39800\,
            I => \N__39706\
        );

    \I__8645\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39693\
        );

    \I__8644\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39693\
        );

    \I__8643\ : InMux
    port map (
            O => \N__39795\,
            I => \N__39693\
        );

    \I__8642\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39693\
        );

    \I__8641\ : InMux
    port map (
            O => \N__39791\,
            I => \N__39693\
        );

    \I__8640\ : InMux
    port map (
            O => \N__39788\,
            I => \N__39693\
        );

    \I__8639\ : InMux
    port map (
            O => \N__39787\,
            I => \N__39686\
        );

    \I__8638\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39686\
        );

    \I__8637\ : InMux
    port map (
            O => \N__39785\,
            I => \N__39686\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__39782\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__39779\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__39768\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8633\ : Odrv12
    port map (
            O => \N__39765\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__39758\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__39747\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__39730\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__39713\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__39706\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8627\ : LocalMux
    port map (
            O => \N__39693\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__39686\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__8625\ : CascadeMux
    port map (
            O => \N__39663\,
            I => \N__39660\
        );

    \I__8624\ : InMux
    port map (
            O => \N__39660\,
            I => \N__39657\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__39657\,
            I => \N__39654\
        );

    \I__8622\ : Span4Mux_v
    port map (
            O => \N__39654\,
            I => \N__39651\
        );

    \I__8621\ : Span4Mux_h
    port map (
            O => \N__39651\,
            I => \N__39648\
        );

    \I__8620\ : Odrv4
    port map (
            O => \N__39648\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__8619\ : InMux
    port map (
            O => \N__39645\,
            I => \N__39642\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__39642\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__8617\ : InMux
    port map (
            O => \N__39639\,
            I => \N__39636\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39633\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__39633\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__8614\ : InMux
    port map (
            O => \N__39630\,
            I => \N__39627\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__39627\,
            I => \N__39624\
        );

    \I__8612\ : Odrv4
    port map (
            O => \N__39624\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__8611\ : InMux
    port map (
            O => \N__39621\,
            I => \N__39618\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__39618\,
            I => \N__39615\
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__39615\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__8608\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39609\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__39609\,
            I => \N__39606\
        );

    \I__8606\ : Odrv4
    port map (
            O => \N__39606\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__8605\ : InMux
    port map (
            O => \N__39603\,
            I => \N__39600\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__39600\,
            I => \N__39596\
        );

    \I__8603\ : InMux
    port map (
            O => \N__39599\,
            I => \N__39593\
        );

    \I__8602\ : Span4Mux_h
    port map (
            O => \N__39596\,
            I => \N__39590\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__39593\,
            I => \N__39587\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__39590\,
            I => \N__39584\
        );

    \I__8599\ : Span4Mux_v
    port map (
            O => \N__39587\,
            I => \N__39580\
        );

    \I__8598\ : Span4Mux_v
    port map (
            O => \N__39584\,
            I => \N__39577\
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__39583\,
            I => \N__39572\
        );

    \I__8596\ : Span4Mux_v
    port map (
            O => \N__39580\,
            I => \N__39569\
        );

    \I__8595\ : Span4Mux_v
    port map (
            O => \N__39577\,
            I => \N__39566\
        );

    \I__8594\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39563\
        );

    \I__8593\ : InMux
    port map (
            O => \N__39575\,
            I => \N__39560\
        );

    \I__8592\ : InMux
    port map (
            O => \N__39572\,
            I => \N__39557\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__39569\,
            I => \N__39554\
        );

    \I__8590\ : Span4Mux_v
    port map (
            O => \N__39566\,
            I => \N__39551\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__39563\,
            I => \N__39548\
        );

    \I__8588\ : LocalMux
    port map (
            O => \N__39560\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__39557\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8586\ : Odrv4
    port map (
            O => \N__39554\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8585\ : Odrv4
    port map (
            O => \N__39551\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8584\ : Odrv4
    port map (
            O => \N__39548\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__8583\ : IoInMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__39534\,
            I => \N__39531\
        );

    \I__8581\ : Span12Mux_s1_v
    port map (
            O => \N__39531\,
            I => \N__39528\
        );

    \I__8580\ : Span12Mux_v
    port map (
            O => \N__39528\,
            I => \N__39524\
        );

    \I__8579\ : InMux
    port map (
            O => \N__39527\,
            I => \N__39521\
        );

    \I__8578\ : Odrv12
    port map (
            O => \N__39524\,
            I => \T01_c\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__39521\,
            I => \T01_c\
        );

    \I__8576\ : InMux
    port map (
            O => \N__39516\,
            I => \N__39513\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__39513\,
            I => \N__39510\
        );

    \I__8574\ : Odrv4
    port map (
            O => \N__39510\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__8573\ : InMux
    port map (
            O => \N__39507\,
            I => \N__39504\
        );

    \I__8572\ : LocalMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__8571\ : Odrv4
    port map (
            O => \N__39501\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__8570\ : InMux
    port map (
            O => \N__39498\,
            I => \N__39494\
        );

    \I__8569\ : InMux
    port map (
            O => \N__39497\,
            I => \N__39491\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__39494\,
            I => \N__39487\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__39491\,
            I => \N__39484\
        );

    \I__8566\ : InMux
    port map (
            O => \N__39490\,
            I => \N__39481\
        );

    \I__8565\ : Span4Mux_h
    port map (
            O => \N__39487\,
            I => \N__39477\
        );

    \I__8564\ : Span4Mux_h
    port map (
            O => \N__39484\,
            I => \N__39472\
        );

    \I__8563\ : LocalMux
    port map (
            O => \N__39481\,
            I => \N__39472\
        );

    \I__8562\ : InMux
    port map (
            O => \N__39480\,
            I => \N__39469\
        );

    \I__8561\ : Odrv4
    port map (
            O => \N__39477\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8560\ : Odrv4
    port map (
            O => \N__39472\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8559\ : LocalMux
    port map (
            O => \N__39469\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__8558\ : InMux
    port map (
            O => \N__39462\,
            I => \N__39459\
        );

    \I__8557\ : LocalMux
    port map (
            O => \N__39459\,
            I => \N__39456\
        );

    \I__8556\ : Odrv4
    port map (
            O => \N__39456\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__8555\ : InMux
    port map (
            O => \N__39453\,
            I => \N__39449\
        );

    \I__8554\ : CascadeMux
    port map (
            O => \N__39452\,
            I => \N__39446\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39441\
        );

    \I__8552\ : InMux
    port map (
            O => \N__39446\,
            I => \N__39438\
        );

    \I__8551\ : InMux
    port map (
            O => \N__39445\,
            I => \N__39432\
        );

    \I__8550\ : InMux
    port map (
            O => \N__39444\,
            I => \N__39432\
        );

    \I__8549\ : Span4Mux_v
    port map (
            O => \N__39441\,
            I => \N__39429\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__39438\,
            I => \N__39426\
        );

    \I__8547\ : InMux
    port map (
            O => \N__39437\,
            I => \N__39423\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__39432\,
            I => \N__39420\
        );

    \I__8545\ : Odrv4
    port map (
            O => \N__39429\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8544\ : Odrv12
    port map (
            O => \N__39426\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8543\ : LocalMux
    port map (
            O => \N__39423\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8542\ : Odrv4
    port map (
            O => \N__39420\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__8541\ : InMux
    port map (
            O => \N__39411\,
            I => \N__39408\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__39408\,
            I => \N__39403\
        );

    \I__8539\ : InMux
    port map (
            O => \N__39407\,
            I => \N__39400\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39406\,
            I => \N__39397\
        );

    \I__8537\ : Span4Mux_v
    port map (
            O => \N__39403\,
            I => \N__39394\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__39400\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8535\ : LocalMux
    port map (
            O => \N__39397\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8534\ : Odrv4
    port map (
            O => \N__39394\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__8533\ : CascadeMux
    port map (
            O => \N__39387\,
            I => \N__39384\
        );

    \I__8532\ : InMux
    port map (
            O => \N__39384\,
            I => \N__39381\
        );

    \I__8531\ : LocalMux
    port map (
            O => \N__39381\,
            I => \N__39378\
        );

    \I__8530\ : Span4Mux_v
    port map (
            O => \N__39378\,
            I => \N__39375\
        );

    \I__8529\ : Span4Mux_h
    port map (
            O => \N__39375\,
            I => \N__39372\
        );

    \I__8528\ : Odrv4
    port map (
            O => \N__39372\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__8527\ : InMux
    port map (
            O => \N__39369\,
            I => \N__39366\
        );

    \I__8526\ : LocalMux
    port map (
            O => \N__39366\,
            I => \N__39361\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39365\,
            I => \N__39358\
        );

    \I__8524\ : InMux
    port map (
            O => \N__39364\,
            I => \N__39355\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__39361\,
            I => \N__39350\
        );

    \I__8522\ : LocalMux
    port map (
            O => \N__39358\,
            I => \N__39350\
        );

    \I__8521\ : LocalMux
    port map (
            O => \N__39355\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__39350\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__8519\ : CascadeMux
    port map (
            O => \N__39345\,
            I => \N__39342\
        );

    \I__8518\ : InMux
    port map (
            O => \N__39342\,
            I => \N__39339\
        );

    \I__8517\ : LocalMux
    port map (
            O => \N__39339\,
            I => \N__39336\
        );

    \I__8516\ : Sp12to4
    port map (
            O => \N__39336\,
            I => \N__39333\
        );

    \I__8515\ : Span12Mux_v
    port map (
            O => \N__39333\,
            I => \N__39330\
        );

    \I__8514\ : Odrv12
    port map (
            O => \N__39330\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__8513\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39324\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39324\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39321\,
            I => \N__39318\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__39318\,
            I => \N__39315\
        );

    \I__8509\ : Odrv4
    port map (
            O => \N__39315\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__8508\ : InMux
    port map (
            O => \N__39312\,
            I => \N__39309\
        );

    \I__8507\ : LocalMux
    port map (
            O => \N__39309\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39306\,
            I => \N__39303\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__39303\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__8504\ : InMux
    port map (
            O => \N__39300\,
            I => \N__39297\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__39297\,
            I => \N__39294\
        );

    \I__8502\ : Odrv4
    port map (
            O => \N__39294\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__8501\ : InMux
    port map (
            O => \N__39291\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__8500\ : InMux
    port map (
            O => \N__39288\,
            I => \bfn_16_14_0_\
        );

    \I__8499\ : InMux
    port map (
            O => \N__39285\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__8498\ : InMux
    port map (
            O => \N__39282\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__8497\ : InMux
    port map (
            O => \N__39279\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__8496\ : InMux
    port map (
            O => \N__39276\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__8495\ : CascadeMux
    port map (
            O => \N__39273\,
            I => \N__39268\
        );

    \I__8494\ : CascadeMux
    port map (
            O => \N__39272\,
            I => \N__39265\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39271\,
            I => \N__39258\
        );

    \I__8492\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39258\
        );

    \I__8491\ : InMux
    port map (
            O => \N__39265\,
            I => \N__39258\
        );

    \I__8490\ : LocalMux
    port map (
            O => \N__39258\,
            I => \N__39254\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39257\,
            I => \N__39251\
        );

    \I__8488\ : Span4Mux_h
    port map (
            O => \N__39254\,
            I => \N__39248\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__39251\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__39248\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39243\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39240\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__8483\ : CascadeMux
    port map (
            O => \N__39237\,
            I => \N__39234\
        );

    \I__8482\ : InMux
    port map (
            O => \N__39234\,
            I => \N__39225\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39233\,
            I => \N__39225\
        );

    \I__8480\ : InMux
    port map (
            O => \N__39232\,
            I => \N__39225\
        );

    \I__8479\ : LocalMux
    port map (
            O => \N__39225\,
            I => \N__39221\
        );

    \I__8478\ : InMux
    port map (
            O => \N__39224\,
            I => \N__39218\
        );

    \I__8477\ : Span4Mux_v
    port map (
            O => \N__39221\,
            I => \N__39215\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39218\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8475\ : Odrv4
    port map (
            O => \N__39215\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__8474\ : InMux
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__39207\,
            I => \N__39203\
        );

    \I__8472\ : InMux
    port map (
            O => \N__39206\,
            I => \N__39200\
        );

    \I__8471\ : Span4Mux_h
    port map (
            O => \N__39203\,
            I => \N__39197\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__39200\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8469\ : Odrv4
    port map (
            O => \N__39197\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__8468\ : InMux
    port map (
            O => \N__39192\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__8467\ : CascadeMux
    port map (
            O => \N__39189\,
            I => \N__39186\
        );

    \I__8466\ : InMux
    port map (
            O => \N__39186\,
            I => \N__39179\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39185\,
            I => \N__39179\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39184\,
            I => \N__39176\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__39179\,
            I => \N__39173\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__39176\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8461\ : Odrv4
    port map (
            O => \N__39173\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__8460\ : InMux
    port map (
            O => \N__39168\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__8459\ : InMux
    port map (
            O => \N__39165\,
            I => \N__39158\
        );

    \I__8458\ : InMux
    port map (
            O => \N__39164\,
            I => \N__39158\
        );

    \I__8457\ : InMux
    port map (
            O => \N__39163\,
            I => \N__39155\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__39158\,
            I => \N__39152\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__39155\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8454\ : Odrv4
    port map (
            O => \N__39152\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39147\,
            I => \bfn_16_13_0_\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39144\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39141\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__39138\,
            I => \N__39134\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39137\,
            I => \N__39128\
        );

    \I__8448\ : InMux
    port map (
            O => \N__39134\,
            I => \N__39128\
        );

    \I__8447\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39125\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__39128\,
            I => \N__39122\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39125\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8444\ : Odrv4
    port map (
            O => \N__39122\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__8443\ : InMux
    port map (
            O => \N__39117\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__8442\ : InMux
    port map (
            O => \N__39114\,
            I => \N__39107\
        );

    \I__8441\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39107\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39112\,
            I => \N__39104\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__39107\,
            I => \N__39101\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__39104\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8437\ : Odrv4
    port map (
            O => \N__39101\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__8436\ : InMux
    port map (
            O => \N__39096\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__8435\ : CascadeMux
    port map (
            O => \N__39093\,
            I => \N__39090\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39090\,
            I => \N__39084\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39089\,
            I => \N__39084\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__39084\,
            I => \N__39080\
        );

    \I__8431\ : InMux
    port map (
            O => \N__39083\,
            I => \N__39077\
        );

    \I__8430\ : Span4Mux_h
    port map (
            O => \N__39080\,
            I => \N__39074\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__39077\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8428\ : Odrv4
    port map (
            O => \N__39074\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__8427\ : InMux
    port map (
            O => \N__39069\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39066\,
            I => \N__39060\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39065\,
            I => \N__39060\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__39060\,
            I => \N__39056\
        );

    \I__8423\ : InMux
    port map (
            O => \N__39059\,
            I => \N__39053\
        );

    \I__8422\ : Span4Mux_h
    port map (
            O => \N__39056\,
            I => \N__39050\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__39053\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__39050\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__8419\ : InMux
    port map (
            O => \N__39045\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__8418\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39038\
        );

    \I__8417\ : InMux
    port map (
            O => \N__39041\,
            I => \N__39035\
        );

    \I__8416\ : LocalMux
    port map (
            O => \N__39038\,
            I => \N__39032\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__39035\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8414\ : Odrv4
    port map (
            O => \N__39032\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39027\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39024\,
            I => \N__39020\
        );

    \I__8411\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39017\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__39020\,
            I => \N__39014\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__39017\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8408\ : Odrv4
    port map (
            O => \N__39014\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__8407\ : InMux
    port map (
            O => \N__39009\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__8406\ : InMux
    port map (
            O => \N__39006\,
            I => \N__39002\
        );

    \I__8405\ : InMux
    port map (
            O => \N__39005\,
            I => \N__38999\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__39002\,
            I => \N__38996\
        );

    \I__8403\ : LocalMux
    port map (
            O => \N__38999\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8402\ : Odrv4
    port map (
            O => \N__38996\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__8401\ : InMux
    port map (
            O => \N__38991\,
            I => \bfn_16_12_0_\
        );

    \I__8400\ : InMux
    port map (
            O => \N__38988\,
            I => \N__38984\
        );

    \I__8399\ : InMux
    port map (
            O => \N__38987\,
            I => \N__38981\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__38984\,
            I => \N__38978\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__38981\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8396\ : Odrv4
    port map (
            O => \N__38978\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__8395\ : InMux
    port map (
            O => \N__38973\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__8394\ : InMux
    port map (
            O => \N__38970\,
            I => \N__38966\
        );

    \I__8393\ : InMux
    port map (
            O => \N__38969\,
            I => \N__38963\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__38966\,
            I => \N__38960\
        );

    \I__8391\ : LocalMux
    port map (
            O => \N__38963\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8390\ : Odrv4
    port map (
            O => \N__38960\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__8389\ : InMux
    port map (
            O => \N__38955\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__8388\ : InMux
    port map (
            O => \N__38952\,
            I => \N__38948\
        );

    \I__8387\ : InMux
    port map (
            O => \N__38951\,
            I => \N__38945\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__38948\,
            I => \N__38942\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__38945\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8384\ : Odrv4
    port map (
            O => \N__38942\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__8383\ : InMux
    port map (
            O => \N__38937\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__8382\ : InMux
    port map (
            O => \N__38934\,
            I => \N__38930\
        );

    \I__8381\ : InMux
    port map (
            O => \N__38933\,
            I => \N__38927\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__38930\,
            I => \N__38924\
        );

    \I__8379\ : LocalMux
    port map (
            O => \N__38927\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__38924\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__8377\ : InMux
    port map (
            O => \N__38919\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__8376\ : InMux
    port map (
            O => \N__38916\,
            I => \N__38912\
        );

    \I__8375\ : InMux
    port map (
            O => \N__38915\,
            I => \N__38909\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__38912\,
            I => \N__38906\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__38909\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8372\ : Odrv12
    port map (
            O => \N__38906\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__8371\ : InMux
    port map (
            O => \N__38901\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__8370\ : InMux
    port map (
            O => \N__38898\,
            I => \N__38895\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__38895\,
            I => \N__38892\
        );

    \I__8368\ : Odrv12
    port map (
            O => \N__38892\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__8367\ : InMux
    port map (
            O => \N__38889\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_28\
        );

    \I__8366\ : InMux
    port map (
            O => \N__38886\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__8365\ : InMux
    port map (
            O => \N__38883\,
            I => \N__38877\
        );

    \I__8364\ : InMux
    port map (
            O => \N__38882\,
            I => \N__38877\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__8362\ : Span4Mux_v
    port map (
            O => \N__38874\,
            I => \N__38871\
        );

    \I__8361\ : Odrv4
    port map (
            O => \N__38871\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__8360\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38865\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__38865\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__8358\ : CascadeMux
    port map (
            O => \N__38862\,
            I => \N__38859\
        );

    \I__8357\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38856\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__38856\,
            I => \N__38851\
        );

    \I__8355\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38848\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__38854\,
            I => \N__38845\
        );

    \I__8353\ : Span4Mux_v
    port map (
            O => \N__38851\,
            I => \N__38842\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__38848\,
            I => \N__38839\
        );

    \I__8351\ : InMux
    port map (
            O => \N__38845\,
            I => \N__38836\
        );

    \I__8350\ : Span4Mux_h
    port map (
            O => \N__38842\,
            I => \N__38833\
        );

    \I__8349\ : Span4Mux_v
    port map (
            O => \N__38839\,
            I => \N__38830\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__38836\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8347\ : Odrv4
    port map (
            O => \N__38833\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8346\ : Odrv4
    port map (
            O => \N__38830\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__8345\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38819\
        );

    \I__8344\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38816\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__38819\,
            I => \N__38813\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__38816\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8341\ : Odrv4
    port map (
            O => \N__38813\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__8340\ : InMux
    port map (
            O => \N__38808\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__8339\ : CascadeMux
    port map (
            O => \N__38805\,
            I => \N__38802\
        );

    \I__8338\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38799\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__38799\,
            I => \N__38796\
        );

    \I__8336\ : Odrv4
    port map (
            O => \N__38796\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\
        );

    \I__8335\ : InMux
    port map (
            O => \N__38793\,
            I => \N__38790\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__38790\,
            I => \N__38786\
        );

    \I__8333\ : InMux
    port map (
            O => \N__38789\,
            I => \N__38783\
        );

    \I__8332\ : Span4Mux_h
    port map (
            O => \N__38786\,
            I => \N__38780\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__38783\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8330\ : Odrv4
    port map (
            O => \N__38780\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__8329\ : InMux
    port map (
            O => \N__38775\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__8328\ : InMux
    port map (
            O => \N__38772\,
            I => \N__38768\
        );

    \I__8327\ : InMux
    port map (
            O => \N__38771\,
            I => \N__38765\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__38768\,
            I => \N__38762\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__38765\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8324\ : Odrv12
    port map (
            O => \N__38762\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__8323\ : InMux
    port map (
            O => \N__38757\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__8322\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38750\
        );

    \I__8321\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38747\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__38750\,
            I => \N__38744\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__38747\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8318\ : Odrv4
    port map (
            O => \N__38744\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__8317\ : InMux
    port map (
            O => \N__38739\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__8316\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__38733\,
            I => \N__38729\
        );

    \I__8314\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38726\
        );

    \I__8313\ : Span4Mux_h
    port map (
            O => \N__38729\,
            I => \N__38723\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__38726\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8311\ : Odrv4
    port map (
            O => \N__38723\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__8310\ : InMux
    port map (
            O => \N__38718\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__8309\ : CascadeMux
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__8308\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38709\
        );

    \I__8307\ : LocalMux
    port map (
            O => \N__38709\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__8306\ : CascadeMux
    port map (
            O => \N__38706\,
            I => \N__38703\
        );

    \I__8305\ : InMux
    port map (
            O => \N__38703\,
            I => \N__38700\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__38700\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__8303\ : InMux
    port map (
            O => \N__38697\,
            I => \N__38694\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__38694\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__8301\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38688\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__38688\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__8299\ : CascadeMux
    port map (
            O => \N__38685\,
            I => \N__38682\
        );

    \I__8298\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38679\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__38679\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__8296\ : InMux
    port map (
            O => \N__38676\,
            I => \N__38673\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__38673\,
            I => \N__38670\
        );

    \I__8294\ : Odrv12
    port map (
            O => \N__38670\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__8293\ : CascadeMux
    port map (
            O => \N__38667\,
            I => \N__38664\
        );

    \I__8292\ : InMux
    port map (
            O => \N__38664\,
            I => \N__38661\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__38661\,
            I => \N__38658\
        );

    \I__8290\ : Span4Mux_v
    port map (
            O => \N__38658\,
            I => \N__38655\
        );

    \I__8289\ : Odrv4
    port map (
            O => \N__38655\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__8288\ : InMux
    port map (
            O => \N__38652\,
            I => \N__38649\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__38649\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__8286\ : CascadeMux
    port map (
            O => \N__38646\,
            I => \N__38643\
        );

    \I__8285\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38640\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__38640\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__8283\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38634\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__38634\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__8281\ : CascadeMux
    port map (
            O => \N__38631\,
            I => \N__38628\
        );

    \I__8280\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38625\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__38625\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__8278\ : InMux
    port map (
            O => \N__38622\,
            I => \N__38619\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__38619\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__8276\ : CascadeMux
    port map (
            O => \N__38616\,
            I => \N__38613\
        );

    \I__8275\ : InMux
    port map (
            O => \N__38613\,
            I => \N__38610\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__38610\,
            I => \N__38607\
        );

    \I__8273\ : Odrv4
    port map (
            O => \N__38607\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__8272\ : CascadeMux
    port map (
            O => \N__38604\,
            I => \N__38601\
        );

    \I__8271\ : InMux
    port map (
            O => \N__38601\,
            I => \N__38598\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__38598\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__8269\ : InMux
    port map (
            O => \N__38595\,
            I => \N__38592\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__38592\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__8267\ : CascadeMux
    port map (
            O => \N__38589\,
            I => \N__38586\
        );

    \I__8266\ : InMux
    port map (
            O => \N__38586\,
            I => \N__38583\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__38583\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__8264\ : InMux
    port map (
            O => \N__38580\,
            I => \N__38577\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__38577\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__38574\,
            I => \N__38571\
        );

    \I__8261\ : InMux
    port map (
            O => \N__38571\,
            I => \N__38568\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__38568\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__8259\ : InMux
    port map (
            O => \N__38565\,
            I => \N__38562\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__38562\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__8257\ : CascadeMux
    port map (
            O => \N__38559\,
            I => \N__38556\
        );

    \I__8256\ : InMux
    port map (
            O => \N__38556\,
            I => \N__38553\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__38553\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__8254\ : CascadeMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__8253\ : InMux
    port map (
            O => \N__38547\,
            I => \N__38544\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__38544\,
            I => \N__38541\
        );

    \I__8251\ : Odrv4
    port map (
            O => \N__38541\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__8250\ : InMux
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__38535\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__38532\,
            I => \N__38529\
        );

    \I__8247\ : InMux
    port map (
            O => \N__38529\,
            I => \N__38526\
        );

    \I__8246\ : LocalMux
    port map (
            O => \N__38526\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__8245\ : InMux
    port map (
            O => \N__38523\,
            I => \N__38520\
        );

    \I__8244\ : LocalMux
    port map (
            O => \N__38520\,
            I => \N__38517\
        );

    \I__8243\ : Odrv4
    port map (
            O => \N__38517\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__8242\ : CascadeMux
    port map (
            O => \N__38514\,
            I => \N__38511\
        );

    \I__8241\ : InMux
    port map (
            O => \N__38511\,
            I => \N__38508\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__38508\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__8239\ : InMux
    port map (
            O => \N__38505\,
            I => \N__38502\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__38502\,
            I => \N__38499\
        );

    \I__8237\ : Odrv12
    port map (
            O => \N__38499\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__8236\ : CascadeMux
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__8235\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__38490\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__8233\ : InMux
    port map (
            O => \N__38487\,
            I => \N__38484\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__38484\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__8231\ : CascadeMux
    port map (
            O => \N__38481\,
            I => \N__38478\
        );

    \I__8230\ : InMux
    port map (
            O => \N__38478\,
            I => \N__38475\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__38475\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__38472\,
            I => \N__38469\
        );

    \I__8227\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38466\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__38466\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__8225\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38460\
        );

    \I__8224\ : LocalMux
    port map (
            O => \N__38460\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__8223\ : CascadeMux
    port map (
            O => \N__38457\,
            I => \N__38452\
        );

    \I__8222\ : CascadeMux
    port map (
            O => \N__38456\,
            I => \N__38449\
        );

    \I__8221\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38443\
        );

    \I__8220\ : InMux
    port map (
            O => \N__38452\,
            I => \N__38443\
        );

    \I__8219\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38438\
        );

    \I__8218\ : InMux
    port map (
            O => \N__38448\,
            I => \N__38438\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__38443\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__38438\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__8215\ : IoInMux
    port map (
            O => \N__38433\,
            I => \N__38430\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__38430\,
            I => \N__38427\
        );

    \I__8213\ : IoSpan4Mux
    port map (
            O => \N__38427\,
            I => \N__38424\
        );

    \I__8212\ : Sp12to4
    port map (
            O => \N__38424\,
            I => \N__38421\
        );

    \I__8211\ : Span12Mux_s6_v
    port map (
            O => \N__38421\,
            I => \N__38418\
        );

    \I__8210\ : Span12Mux_v
    port map (
            O => \N__38418\,
            I => \N__38414\
        );

    \I__8209\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38411\
        );

    \I__8208\ : Odrv12
    port map (
            O => \N__38414\,
            I => \T12_c\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__38411\,
            I => \T12_c\
        );

    \I__8206\ : CascadeMux
    port map (
            O => \N__38406\,
            I => \N__38403\
        );

    \I__8205\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38399\
        );

    \I__8204\ : InMux
    port map (
            O => \N__38402\,
            I => \N__38396\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__38399\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__38396\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__38391\,
            I => \N__38387\
        );

    \I__8200\ : InMux
    port map (
            O => \N__38390\,
            I => \N__38380\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38380\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38386\,
            I => \N__38377\
        );

    \I__8197\ : InMux
    port map (
            O => \N__38385\,
            I => \N__38374\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__38380\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__38377\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38374\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__8193\ : CascadeMux
    port map (
            O => \N__38367\,
            I => \N__38363\
        );

    \I__8192\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38355\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38363\,
            I => \N__38355\
        );

    \I__8190\ : InMux
    port map (
            O => \N__38362\,
            I => \N__38352\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38361\,
            I => \N__38347\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38360\,
            I => \N__38347\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__38355\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__38352\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38347\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__8184\ : CascadeMux
    port map (
            O => \N__38340\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38337\,
            I => \N__38331\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38336\,
            I => \N__38331\
        );

    \I__8181\ : LocalMux
    port map (
            O => \N__38331\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__38328\,
            I => \N__38325\
        );

    \I__8179\ : InMux
    port map (
            O => \N__38325\,
            I => \N__38319\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38324\,
            I => \N__38319\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__38319\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__8176\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38311\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38308\
        );

    \I__8174\ : InMux
    port map (
            O => \N__38314\,
            I => \N__38305\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__38311\,
            I => \N__38302\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38308\,
            I => \N__38299\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__38305\,
            I => \N__38296\
        );

    \I__8170\ : Odrv12
    port map (
            O => \N__38302\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8169\ : Odrv12
    port map (
            O => \N__38299\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__38296\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38289\,
            I => \N__38286\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38286\,
            I => \N__38283\
        );

    \I__8165\ : Odrv12
    port map (
            O => \N__38283\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__38280\,
            I => \N__38277\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38271\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38271\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38271\,
            I => \N__38267\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38270\,
            I => \N__38264\
        );

    \I__8159\ : Span4Mux_h
    port map (
            O => \N__38267\,
            I => \N__38261\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__38264\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__38261\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__8156\ : InMux
    port map (
            O => \N__38256\,
            I => \N__38252\
        );

    \I__8155\ : InMux
    port map (
            O => \N__38255\,
            I => \N__38249\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38252\,
            I => \N__38242\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38249\,
            I => \N__38242\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38248\,
            I => \N__38239\
        );

    \I__8151\ : InMux
    port map (
            O => \N__38247\,
            I => \N__38236\
        );

    \I__8150\ : Span4Mux_h
    port map (
            O => \N__38242\,
            I => \N__38233\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__38239\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__38236\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__8147\ : Odrv4
    port map (
            O => \N__38233\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__8146\ : ClkMux
    port map (
            O => \N__38226\,
            I => \N__38220\
        );

    \I__8145\ : ClkMux
    port map (
            O => \N__38225\,
            I => \N__38220\
        );

    \I__8144\ : GlobalMux
    port map (
            O => \N__38220\,
            I => \N__38217\
        );

    \I__8143\ : gio2CtrlBuf
    port map (
            O => \N__38217\,
            I => delay_tr_input_c_g
        );

    \I__8142\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38207\
        );

    \I__8141\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38207\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38204\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__38207\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__38204\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__8137\ : InMux
    port map (
            O => \N__38199\,
            I => \N__38195\
        );

    \I__8136\ : InMux
    port map (
            O => \N__38198\,
            I => \N__38192\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__38195\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__38192\,
            I => \phase_controller_inst2.state_RNI9M3OZ0Z_0\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38187\,
            I => \N__38184\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__38184\,
            I => \phase_controller_inst2.start_timer_tr_RNO_0_0\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38181\,
            I => \N__38177\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38180\,
            I => \N__38174\
        );

    \I__8129\ : LocalMux
    port map (
            O => \N__38177\,
            I => \N__38170\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__38174\,
            I => \N__38167\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38173\,
            I => \N__38164\
        );

    \I__8126\ : Span4Mux_h
    port map (
            O => \N__38170\,
            I => \N__38161\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__38167\,
            I => \N__38158\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__38164\,
            I => \N__38155\
        );

    \I__8123\ : Span4Mux_h
    port map (
            O => \N__38161\,
            I => \N__38152\
        );

    \I__8122\ : Span4Mux_h
    port map (
            O => \N__38158\,
            I => \N__38149\
        );

    \I__8121\ : Span12Mux_h
    port map (
            O => \N__38155\,
            I => \N__38146\
        );

    \I__8120\ : Span4Mux_h
    port map (
            O => \N__38152\,
            I => \N__38143\
        );

    \I__8119\ : Span4Mux_h
    port map (
            O => \N__38149\,
            I => \N__38140\
        );

    \I__8118\ : Odrv12
    port map (
            O => \N__38146\,
            I => il_max_comp2_c
        );

    \I__8117\ : Odrv4
    port map (
            O => \N__38143\,
            I => il_max_comp2_c
        );

    \I__8116\ : Odrv4
    port map (
            O => \N__38140\,
            I => il_max_comp2_c
        );

    \I__8115\ : InMux
    port map (
            O => \N__38133\,
            I => \N__38128\
        );

    \I__8114\ : InMux
    port map (
            O => \N__38132\,
            I => \N__38123\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38123\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__38128\,
            I => \N__38117\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__38123\,
            I => \N__38117\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38114\
        );

    \I__8109\ : Span4Mux_h
    port map (
            O => \N__38117\,
            I => \N__38111\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__38114\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__8107\ : Odrv4
    port map (
            O => \N__38111\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38106\,
            I => \N__38101\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38105\,
            I => \N__38098\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38104\,
            I => \N__38095\
        );

    \I__8103\ : LocalMux
    port map (
            O => \N__38101\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__8102\ : LocalMux
    port map (
            O => \N__38098\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__38095\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__8100\ : InMux
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__38085\,
            I => \N__38082\
        );

    \I__8098\ : Odrv12
    port map (
            O => \N__38082\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8097\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38076\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38076\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__38073\,
            I => \N__38069\
        );

    \I__8094\ : InMux
    port map (
            O => \N__38072\,
            I => \N__38064\
        );

    \I__8093\ : InMux
    port map (
            O => \N__38069\,
            I => \N__38064\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38064\,
            I => \N__38060\
        );

    \I__8091\ : InMux
    port map (
            O => \N__38063\,
            I => \N__38057\
        );

    \I__8090\ : Span4Mux_v
    port map (
            O => \N__38060\,
            I => \N__38054\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__38057\,
            I => \N__38051\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__38054\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8087\ : Odrv4
    port map (
            O => \N__38051\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__8086\ : InMux
    port map (
            O => \N__38046\,
            I => \N__38043\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38043\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8084\ : InMux
    port map (
            O => \N__38040\,
            I => \N__38019\
        );

    \I__8083\ : InMux
    port map (
            O => \N__38039\,
            I => \N__38019\
        );

    \I__8082\ : InMux
    port map (
            O => \N__38038\,
            I => \N__38019\
        );

    \I__8081\ : InMux
    port map (
            O => \N__38037\,
            I => \N__38019\
        );

    \I__8080\ : InMux
    port map (
            O => \N__38036\,
            I => \N__38019\
        );

    \I__8079\ : InMux
    port map (
            O => \N__38035\,
            I => \N__38019\
        );

    \I__8078\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38019\
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__38019\,
            I => \N__37999\
        );

    \I__8076\ : InMux
    port map (
            O => \N__38018\,
            I => \N__37994\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38017\,
            I => \N__37994\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38016\,
            I => \N__37991\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38015\,
            I => \N__37980\
        );

    \I__8072\ : InMux
    port map (
            O => \N__38014\,
            I => \N__37980\
        );

    \I__8071\ : InMux
    port map (
            O => \N__38013\,
            I => \N__37980\
        );

    \I__8070\ : InMux
    port map (
            O => \N__38012\,
            I => \N__37980\
        );

    \I__8069\ : InMux
    port map (
            O => \N__38011\,
            I => \N__37980\
        );

    \I__8068\ : InMux
    port map (
            O => \N__38010\,
            I => \N__37971\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38009\,
            I => \N__37971\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38008\,
            I => \N__37971\
        );

    \I__8065\ : InMux
    port map (
            O => \N__38007\,
            I => \N__37971\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38006\,
            I => \N__37968\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38005\,
            I => \N__37965\
        );

    \I__8062\ : InMux
    port map (
            O => \N__38004\,
            I => \N__37958\
        );

    \I__8061\ : InMux
    port map (
            O => \N__38003\,
            I => \N__37958\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38002\,
            I => \N__37958\
        );

    \I__8059\ : Span4Mux_v
    port map (
            O => \N__37999\,
            I => \N__37952\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__37994\,
            I => \N__37952\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__37991\,
            I => \N__37947\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__37980\,
            I => \N__37947\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__37971\,
            I => \N__37938\
        );

    \I__8054\ : LocalMux
    port map (
            O => \N__37968\,
            I => \N__37938\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__37965\,
            I => \N__37938\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__37958\,
            I => \N__37938\
        );

    \I__8051\ : InMux
    port map (
            O => \N__37957\,
            I => \N__37935\
        );

    \I__8050\ : Span4Mux_h
    port map (
            O => \N__37952\,
            I => \N__37932\
        );

    \I__8049\ : Span4Mux_h
    port map (
            O => \N__37947\,
            I => \N__37929\
        );

    \I__8048\ : Span4Mux_v
    port map (
            O => \N__37938\,
            I => \N__37926\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__37935\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__37932\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8045\ : Odrv4
    port map (
            O => \N__37929\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8044\ : Odrv4
    port map (
            O => \N__37926\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__8043\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37912\
        );

    \I__8042\ : InMux
    port map (
            O => \N__37916\,
            I => \N__37909\
        );

    \I__8041\ : InMux
    port map (
            O => \N__37915\,
            I => \N__37906\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__37912\,
            I => \N__37901\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__37909\,
            I => \N__37901\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__37906\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8037\ : Odrv12
    port map (
            O => \N__37901\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__8036\ : CascadeMux
    port map (
            O => \N__37896\,
            I => \N__37893\
        );

    \I__8035\ : InMux
    port map (
            O => \N__37893\,
            I => \N__37890\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__37890\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__8033\ : InMux
    port map (
            O => \N__37887\,
            I => \N__37884\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__37884\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__8031\ : CascadeMux
    port map (
            O => \N__37881\,
            I => \N__37878\
        );

    \I__8030\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37875\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__37875\,
            I => \N__37870\
        );

    \I__8028\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37867\
        );

    \I__8027\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37864\
        );

    \I__8026\ : Span4Mux_h
    port map (
            O => \N__37870\,
            I => \N__37859\
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__37867\,
            I => \N__37859\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__37864\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__37859\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__8022\ : CascadeMux
    port map (
            O => \N__37854\,
            I => \N__37851\
        );

    \I__8021\ : InMux
    port map (
            O => \N__37851\,
            I => \N__37848\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__37848\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__37845\,
            I => \N__37842\
        );

    \I__8018\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37839\
        );

    \I__8017\ : LocalMux
    port map (
            O => \N__37839\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__8016\ : CascadeMux
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__8015\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37830\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__37830\,
            I => \N__37825\
        );

    \I__8013\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37822\
        );

    \I__8012\ : InMux
    port map (
            O => \N__37828\,
            I => \N__37819\
        );

    \I__8011\ : Sp12to4
    port map (
            O => \N__37825\,
            I => \N__37814\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__37822\,
            I => \N__37814\
        );

    \I__8009\ : LocalMux
    port map (
            O => \N__37819\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__8008\ : Odrv12
    port map (
            O => \N__37814\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__8007\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37806\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__37806\,
            I => \N__37803\
        );

    \I__8005\ : Odrv12
    port map (
            O => \N__37803\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__8004\ : CascadeMux
    port map (
            O => \N__37800\,
            I => \N__37797\
        );

    \I__8003\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37794\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__37794\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__8001\ : CascadeMux
    port map (
            O => \N__37791\,
            I => \N__37788\
        );

    \I__8000\ : InMux
    port map (
            O => \N__37788\,
            I => \N__37785\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__37785\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__7998\ : CascadeMux
    port map (
            O => \N__37782\,
            I => \N__37779\
        );

    \I__7997\ : InMux
    port map (
            O => \N__37779\,
            I => \N__37776\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__37776\,
            I => \N__37771\
        );

    \I__7995\ : InMux
    port map (
            O => \N__37775\,
            I => \N__37768\
        );

    \I__7994\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37765\
        );

    \I__7993\ : Span4Mux_v
    port map (
            O => \N__37771\,
            I => \N__37762\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__37768\,
            I => \N__37759\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__37765\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__7990\ : Odrv4
    port map (
            O => \N__37762\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__7989\ : Odrv12
    port map (
            O => \N__37759\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__7988\ : CascadeMux
    port map (
            O => \N__37752\,
            I => \N__37749\
        );

    \I__7987\ : InMux
    port map (
            O => \N__37749\,
            I => \N__37746\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__37746\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__7985\ : CascadeMux
    port map (
            O => \N__37743\,
            I => \N__37738\
        );

    \I__7984\ : InMux
    port map (
            O => \N__37742\,
            I => \N__37735\
        );

    \I__7983\ : InMux
    port map (
            O => \N__37741\,
            I => \N__37730\
        );

    \I__7982\ : InMux
    port map (
            O => \N__37738\,
            I => \N__37730\
        );

    \I__7981\ : LocalMux
    port map (
            O => \N__37735\,
            I => \N__37727\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__37730\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__7979\ : Odrv4
    port map (
            O => \N__37727\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__7978\ : InMux
    port map (
            O => \N__37722\,
            I => \N__37719\
        );

    \I__7977\ : LocalMux
    port map (
            O => \N__37719\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__7976\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37713\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__37713\,
            I => \N__37709\
        );

    \I__7974\ : InMux
    port map (
            O => \N__37712\,
            I => \N__37705\
        );

    \I__7973\ : Span4Mux_v
    port map (
            O => \N__37709\,
            I => \N__37702\
        );

    \I__7972\ : InMux
    port map (
            O => \N__37708\,
            I => \N__37699\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37696\
        );

    \I__7970\ : Odrv4
    port map (
            O => \N__37702\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__37699\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__7968\ : Odrv12
    port map (
            O => \N__37696\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__7967\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37686\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__37686\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__7965\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37678\
        );

    \I__7964\ : InMux
    port map (
            O => \N__37682\,
            I => \N__37675\
        );

    \I__7963\ : InMux
    port map (
            O => \N__37681\,
            I => \N__37672\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__37678\,
            I => \N__37669\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__37675\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__7960\ : LocalMux
    port map (
            O => \N__37672\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__7959\ : Odrv4
    port map (
            O => \N__37669\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__7958\ : InMux
    port map (
            O => \N__37662\,
            I => \N__37659\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__37659\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__37656\,
            I => \N__37651\
        );

    \I__7955\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37648\
        );

    \I__7954\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37645\
        );

    \I__7953\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37642\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__37648\,
            I => \N__37639\
        );

    \I__7951\ : LocalMux
    port map (
            O => \N__37645\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__37642\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__7949\ : Odrv4
    port map (
            O => \N__37639\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__7948\ : CascadeMux
    port map (
            O => \N__37632\,
            I => \N__37629\
        );

    \I__7947\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37626\
        );

    \I__7946\ : LocalMux
    port map (
            O => \N__37626\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__7945\ : CascadeMux
    port map (
            O => \N__37623\,
            I => \N__37620\
        );

    \I__7944\ : InMux
    port map (
            O => \N__37620\,
            I => \N__37617\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__37617\,
            I => \N__37612\
        );

    \I__7942\ : InMux
    port map (
            O => \N__37616\,
            I => \N__37609\
        );

    \I__7941\ : InMux
    port map (
            O => \N__37615\,
            I => \N__37606\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__37612\,
            I => \N__37603\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__37609\,
            I => \N__37600\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__37606\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__7937\ : Odrv4
    port map (
            O => \N__37603\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__7936\ : Odrv12
    port map (
            O => \N__37600\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__7935\ : CascadeMux
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__7934\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37587\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__37587\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__37584\,
            I => \N__37581\
        );

    \I__7931\ : InMux
    port map (
            O => \N__37581\,
            I => \N__37578\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__37578\,
            I => \N__37575\
        );

    \I__7929\ : Span4Mux_h
    port map (
            O => \N__37575\,
            I => \N__37570\
        );

    \I__7928\ : InMux
    port map (
            O => \N__37574\,
            I => \N__37567\
        );

    \I__7927\ : InMux
    port map (
            O => \N__37573\,
            I => \N__37564\
        );

    \I__7926\ : Sp12to4
    port map (
            O => \N__37570\,
            I => \N__37559\
        );

    \I__7925\ : LocalMux
    port map (
            O => \N__37567\,
            I => \N__37559\
        );

    \I__7924\ : LocalMux
    port map (
            O => \N__37564\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__7923\ : Odrv12
    port map (
            O => \N__37559\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__7922\ : InMux
    port map (
            O => \N__37554\,
            I => \N__37551\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__37551\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__7920\ : CascadeMux
    port map (
            O => \N__37548\,
            I => \N__37544\
        );

    \I__7919\ : InMux
    port map (
            O => \N__37547\,
            I => \N__37541\
        );

    \I__7918\ : InMux
    port map (
            O => \N__37544\,
            I => \N__37538\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__37541\,
            I => \N__37532\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__37538\,
            I => \N__37532\
        );

    \I__7915\ : InMux
    port map (
            O => \N__37537\,
            I => \N__37529\
        );

    \I__7914\ : Span4Mux_h
    port map (
            O => \N__37532\,
            I => \N__37526\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__37529\,
            I => \N__37523\
        );

    \I__7912\ : Span4Mux_h
    port map (
            O => \N__37526\,
            I => \N__37518\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__37523\,
            I => \N__37518\
        );

    \I__7910\ : Odrv4
    port map (
            O => \N__37518\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__7909\ : CascadeMux
    port map (
            O => \N__37515\,
            I => \N__37512\
        );

    \I__7908\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37509\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__37509\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__7906\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37503\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__37503\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__37500\,
            I => \N__37495\
        );

    \I__7903\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37492\
        );

    \I__7902\ : InMux
    port map (
            O => \N__37498\,
            I => \N__37487\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37495\,
            I => \N__37487\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37492\,
            I => \N__37484\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__37487\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__37484\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__7897\ : InMux
    port map (
            O => \N__37479\,
            I => \N__37476\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__37476\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37473\,
            I => \N__37468\
        );

    \I__7894\ : InMux
    port map (
            O => \N__37472\,
            I => \N__37465\
        );

    \I__7893\ : InMux
    port map (
            O => \N__37471\,
            I => \N__37462\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__37468\,
            I => \N__37457\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__37465\,
            I => \N__37457\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__37462\,
            I => \N__37454\
        );

    \I__7889\ : Span4Mux_v
    port map (
            O => \N__37457\,
            I => \N__37451\
        );

    \I__7888\ : Span4Mux_v
    port map (
            O => \N__37454\,
            I => \N__37448\
        );

    \I__7887\ : Odrv4
    port map (
            O => \N__37451\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__7886\ : Odrv4
    port map (
            O => \N__37448\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__7885\ : CascadeMux
    port map (
            O => \N__37443\,
            I => \N__37440\
        );

    \I__7884\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37437\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__37437\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__7882\ : InMux
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37431\,
            I => \N__37427\
        );

    \I__7880\ : InMux
    port map (
            O => \N__37430\,
            I => \N__37424\
        );

    \I__7879\ : Span4Mux_h
    port map (
            O => \N__37427\,
            I => \N__37418\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__37424\,
            I => \N__37418\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37423\,
            I => \N__37415\
        );

    \I__7876\ : Span4Mux_v
    port map (
            O => \N__37418\,
            I => \N__37412\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37415\,
            I => \N__37409\
        );

    \I__7874\ : Odrv4
    port map (
            O => \N__37412\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7873\ : Odrv4
    port map (
            O => \N__37409\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__7872\ : CascadeMux
    port map (
            O => \N__37404\,
            I => \N__37401\
        );

    \I__7871\ : InMux
    port map (
            O => \N__37401\,
            I => \N__37398\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__37398\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__7869\ : CascadeMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__7868\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__7866\ : Span4Mux_h
    port map (
            O => \N__37386\,
            I => \N__37383\
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__37383\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__7864\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37376\
        );

    \I__7863\ : InMux
    port map (
            O => \N__37379\,
            I => \N__37373\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__37376\,
            I => \N__37369\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37373\,
            I => \N__37366\
        );

    \I__7860\ : InMux
    port map (
            O => \N__37372\,
            I => \N__37363\
        );

    \I__7859\ : Span4Mux_v
    port map (
            O => \N__37369\,
            I => \N__37360\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__37366\,
            I => \N__37357\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__37363\,
            I => \N__37354\
        );

    \I__7856\ : Odrv4
    port map (
            O => \N__37360\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__37357\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7854\ : Odrv4
    port map (
            O => \N__37354\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__7852\ : InMux
    port map (
            O => \N__37344\,
            I => \N__37341\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__37341\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__7850\ : CascadeMux
    port map (
            O => \N__37338\,
            I => \N__37335\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37332\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__7847\ : Span4Mux_h
    port map (
            O => \N__37329\,
            I => \N__37326\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__37326\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__7845\ : CascadeMux
    port map (
            O => \N__37323\,
            I => \N__37320\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37317\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__37317\,
            I => \N__37314\
        );

    \I__7842\ : Span4Mux_h
    port map (
            O => \N__37314\,
            I => \N__37311\
        );

    \I__7841\ : Odrv4
    port map (
            O => \N__37311\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37308\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37305\,
            I => \bfn_15_16_0_\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37302\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37299\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__7836\ : InMux
    port map (
            O => \N__37296\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37293\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__7834\ : InMux
    port map (
            O => \N__37290\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__37287\,
            I => \N__37284\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37281\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37281\,
            I => \N__37278\
        );

    \I__7830\ : Span4Mux_h
    port map (
            O => \N__37278\,
            I => \N__37275\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__37275\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__37272\,
            I => \N__37269\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37266\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__37266\,
            I => \N__37263\
        );

    \I__7825\ : Span4Mux_h
    port map (
            O => \N__37263\,
            I => \N__37260\
        );

    \I__7824\ : Odrv4
    port map (
            O => \N__37260\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37257\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__7822\ : InMux
    port map (
            O => \N__37254\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__7821\ : InMux
    port map (
            O => \N__37251\,
            I => \bfn_15_15_0_\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37248\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37245\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37242\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__7817\ : CascadeMux
    port map (
            O => \N__37239\,
            I => \N__37236\
        );

    \I__7816\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37229\
        );

    \I__7815\ : InMux
    port map (
            O => \N__37235\,
            I => \N__37229\
        );

    \I__7814\ : InMux
    port map (
            O => \N__37234\,
            I => \N__37226\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__37229\,
            I => \N__37223\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__37226\,
            I => \N__37220\
        );

    \I__7811\ : Span4Mux_v
    port map (
            O => \N__37223\,
            I => \N__37217\
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__37220\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__7809\ : Odrv4
    port map (
            O => \N__37217\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37212\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37209\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37206\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37200\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__37200\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37197\,
            I => \N__37193\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37196\,
            I => \N__37190\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37193\,
            I => \N__37187\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__37190\,
            I => \N__37184\
        );

    \I__7799\ : Span4Mux_v
    port map (
            O => \N__37187\,
            I => \N__37180\
        );

    \I__7798\ : Span4Mux_h
    port map (
            O => \N__37184\,
            I => \N__37177\
        );

    \I__7797\ : InMux
    port map (
            O => \N__37183\,
            I => \N__37174\
        );

    \I__7796\ : Odrv4
    port map (
            O => \N__37180\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7795\ : Odrv4
    port map (
            O => \N__37177\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__37174\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__7793\ : InMux
    port map (
            O => \N__37167\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37164\,
            I => \N__37160\
        );

    \I__7791\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37157\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__37160\,
            I => \N__37152\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37152\
        );

    \I__7788\ : Span4Mux_h
    port map (
            O => \N__37152\,
            I => \N__37148\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37151\,
            I => \N__37145\
        );

    \I__7786\ : Odrv4
    port map (
            O => \N__37148\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__37145\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__7784\ : InMux
    port map (
            O => \N__37140\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__7783\ : InMux
    port map (
            O => \N__37137\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__7782\ : InMux
    port map (
            O => \N__37134\,
            I => \N__37131\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37131\,
            I => \N__37127\
        );

    \I__7780\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37124\
        );

    \I__7779\ : Span4Mux_h
    port map (
            O => \N__37127\,
            I => \N__37119\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__37124\,
            I => \N__37119\
        );

    \I__7777\ : Span4Mux_v
    port map (
            O => \N__37119\,
            I => \N__37115\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37118\,
            I => \N__37112\
        );

    \I__7775\ : Odrv4
    port map (
            O => \N__37115\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37112\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__7773\ : InMux
    port map (
            O => \N__37107\,
            I => \bfn_15_14_0_\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37104\,
            I => \N__37101\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__37101\,
            I => \N__37097\
        );

    \I__7770\ : CascadeMux
    port map (
            O => \N__37100\,
            I => \N__37094\
        );

    \I__7769\ : Span4Mux_v
    port map (
            O => \N__37097\,
            I => \N__37090\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37085\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37085\
        );

    \I__7766\ : Odrv4
    port map (
            O => \N__37090\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__37085\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37080\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37077\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__7762\ : CascadeMux
    port map (
            O => \N__37074\,
            I => \N__37071\
        );

    \I__7761\ : InMux
    port map (
            O => \N__37071\,
            I => \N__37068\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__37068\,
            I => \N__37064\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37067\,
            I => \N__37061\
        );

    \I__7758\ : Span4Mux_h
    port map (
            O => \N__37064\,
            I => \N__37058\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__37061\,
            I => \N__37055\
        );

    \I__7756\ : Span4Mux_v
    port map (
            O => \N__37058\,
            I => \N__37049\
        );

    \I__7755\ : Span4Mux_v
    port map (
            O => \N__37055\,
            I => \N__37049\
        );

    \I__7754\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37046\
        );

    \I__7753\ : Odrv4
    port map (
            O => \N__37049\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37046\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37041\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__37038\,
            I => \N__37035\
        );

    \I__7749\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37031\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__37034\,
            I => \N__37028\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__37031\,
            I => \N__37025\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37022\
        );

    \I__7745\ : Span4Mux_v
    port map (
            O => \N__37025\,
            I => \N__37019\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__37022\,
            I => \N__37016\
        );

    \I__7743\ : Span4Mux_h
    port map (
            O => \N__37019\,
            I => \N__37012\
        );

    \I__7742\ : Span4Mux_h
    port map (
            O => \N__37016\,
            I => \N__37009\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37015\,
            I => \N__37006\
        );

    \I__7740\ : Odrv4
    port map (
            O => \N__37012\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__7739\ : Odrv4
    port map (
            O => \N__37009\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37006\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__7737\ : InMux
    port map (
            O => \N__36999\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__7736\ : InMux
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__36993\,
            I => \N__36990\
        );

    \I__7734\ : Odrv4
    port map (
            O => \N__36990\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__7733\ : InMux
    port map (
            O => \N__36987\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__36984\,
            I => \N__36980\
        );

    \I__7731\ : InMux
    port map (
            O => \N__36983\,
            I => \N__36977\
        );

    \I__7730\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36974\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__36977\,
            I => \N__36971\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__36974\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__7727\ : Odrv4
    port map (
            O => \N__36971\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__7726\ : CascadeMux
    port map (
            O => \N__36966\,
            I => \N__36963\
        );

    \I__7725\ : InMux
    port map (
            O => \N__36963\,
            I => \N__36960\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__36960\,
            I => \N__36957\
        );

    \I__7723\ : Odrv4
    port map (
            O => \N__36957\,
            I => \phase_controller_inst1.stoper_tr.un4_running_df30\
        );

    \I__7722\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__7721\ : LocalMux
    port map (
            O => \N__36951\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\
        );

    \I__7720\ : CascadeMux
    port map (
            O => \N__36948\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__7719\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36942\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__36942\,
            I => \N__36939\
        );

    \I__7717\ : Span4Mux_h
    port map (
            O => \N__36939\,
            I => \N__36936\
        );

    \I__7716\ : Span4Mux_v
    port map (
            O => \N__36936\,
            I => \N__36932\
        );

    \I__7715\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36929\
        );

    \I__7714\ : Odrv4
    port map (
            O => \N__36932\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__36929\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__7712\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36921\
        );

    \I__7711\ : LocalMux
    port map (
            O => \N__36921\,
            I => \N__36917\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__36920\,
            I => \N__36913\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__36917\,
            I => \N__36909\
        );

    \I__7708\ : InMux
    port map (
            O => \N__36916\,
            I => \N__36906\
        );

    \I__7707\ : InMux
    port map (
            O => \N__36913\,
            I => \N__36903\
        );

    \I__7706\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36900\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__36909\,
            I => \N__36897\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__36906\,
            I => \N__36892\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__36903\,
            I => \N__36892\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__36900\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__36897\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7700\ : Odrv4
    port map (
            O => \N__36892\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__7699\ : InMux
    port map (
            O => \N__36885\,
            I => \N__36882\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__36882\,
            I => \N__36878\
        );

    \I__7697\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36875\
        );

    \I__7696\ : Span4Mux_v
    port map (
            O => \N__36878\,
            I => \N__36872\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__36875\,
            I => \N__36869\
        );

    \I__7694\ : Span4Mux_h
    port map (
            O => \N__36872\,
            I => \N__36865\
        );

    \I__7693\ : Span4Mux_v
    port map (
            O => \N__36869\,
            I => \N__36862\
        );

    \I__7692\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36859\
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__36865\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__36862\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__36859\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__7688\ : InMux
    port map (
            O => \N__36852\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__7687\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36844\
        );

    \I__7686\ : InMux
    port map (
            O => \N__36848\,
            I => \N__36841\
        );

    \I__7685\ : InMux
    port map (
            O => \N__36847\,
            I => \N__36838\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__36844\,
            I => \N__36833\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__36841\,
            I => \N__36833\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__36838\,
            I => \N__36830\
        );

    \I__7681\ : Span4Mux_v
    port map (
            O => \N__36833\,
            I => \N__36827\
        );

    \I__7680\ : Span4Mux_h
    port map (
            O => \N__36830\,
            I => \N__36824\
        );

    \I__7679\ : Odrv4
    port map (
            O => \N__36827\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__7678\ : Odrv4
    port map (
            O => \N__36824\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__7677\ : InMux
    port map (
            O => \N__36819\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__7676\ : InMux
    port map (
            O => \N__36816\,
            I => \N__36811\
        );

    \I__7675\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36808\
        );

    \I__7674\ : InMux
    port map (
            O => \N__36814\,
            I => \N__36805\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__36811\,
            I => \N__36802\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__36808\,
            I => \N__36797\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__36805\,
            I => \N__36797\
        );

    \I__7670\ : Span4Mux_h
    port map (
            O => \N__36802\,
            I => \N__36794\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__36797\,
            I => \N__36791\
        );

    \I__7668\ : Odrv4
    port map (
            O => \N__36794\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__7667\ : Odrv4
    port map (
            O => \N__36791\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__7666\ : InMux
    port map (
            O => \N__36786\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__7665\ : InMux
    port map (
            O => \N__36783\,
            I => \N__36780\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__7663\ : Span4Mux_h
    port map (
            O => \N__36777\,
            I => \N__36774\
        );

    \I__7662\ : Span4Mux_h
    port map (
            O => \N__36774\,
            I => \N__36771\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__36771\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__7660\ : InMux
    port map (
            O => \N__36768\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__7659\ : CascadeMux
    port map (
            O => \N__36765\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__7658\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36759\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__36759\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__7656\ : InMux
    port map (
            O => \N__36756\,
            I => \N__36753\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__36753\,
            I => \N__36749\
        );

    \I__7654\ : InMux
    port map (
            O => \N__36752\,
            I => \N__36746\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__36749\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__36746\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__7651\ : CascadeMux
    port map (
            O => \N__36741\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\
        );

    \I__7650\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36730\
        );

    \I__7649\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36730\
        );

    \I__7648\ : InMux
    port map (
            O => \N__36736\,
            I => \N__36727\
        );

    \I__7647\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36724\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__36730\,
            I => \N__36719\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__36727\,
            I => \N__36719\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__36724\,
            I => \N__36716\
        );

    \I__7643\ : Span4Mux_v
    port map (
            O => \N__36719\,
            I => \N__36713\
        );

    \I__7642\ : Odrv4
    port map (
            O => \N__36716\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7641\ : Odrv4
    port map (
            O => \N__36713\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7640\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36705\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__36705\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__7638\ : CascadeMux
    port map (
            O => \N__36702\,
            I => \N__36699\
        );

    \I__7637\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36693\
        );

    \I__7636\ : InMux
    port map (
            O => \N__36698\,
            I => \N__36693\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__36693\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__7634\ : CascadeMux
    port map (
            O => \N__36690\,
            I => \N__36687\
        );

    \I__7633\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36684\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__36684\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__7631\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36678\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__36678\,
            I => \N__36674\
        );

    \I__7629\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36671\
        );

    \I__7628\ : Odrv12
    port map (
            O => \N__36674\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__36671\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__7626\ : CascadeMux
    port map (
            O => \N__36666\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\
        );

    \I__7625\ : InMux
    port map (
            O => \N__36663\,
            I => \N__36658\
        );

    \I__7624\ : InMux
    port map (
            O => \N__36662\,
            I => \N__36653\
        );

    \I__7623\ : InMux
    port map (
            O => \N__36661\,
            I => \N__36653\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__36658\,
            I => \N__36649\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__36653\,
            I => \N__36646\
        );

    \I__7620\ : InMux
    port map (
            O => \N__36652\,
            I => \N__36643\
        );

    \I__7619\ : Sp12to4
    port map (
            O => \N__36649\,
            I => \N__36640\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__36646\,
            I => \N__36637\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__36643\,
            I => \N__36634\
        );

    \I__7616\ : Odrv12
    port map (
            O => \N__36640\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__7615\ : Odrv4
    port map (
            O => \N__36637\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__36634\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__7613\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36621\
        );

    \I__7612\ : InMux
    port map (
            O => \N__36626\,
            I => \N__36621\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__36621\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__7610\ : CascadeMux
    port map (
            O => \N__36618\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\
        );

    \I__7609\ : InMux
    port map (
            O => \N__36615\,
            I => \N__36612\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__36612\,
            I => \N__36608\
        );

    \I__7607\ : InMux
    port map (
            O => \N__36611\,
            I => \N__36605\
        );

    \I__7606\ : Span4Mux_h
    port map (
            O => \N__36608\,
            I => \N__36599\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__36605\,
            I => \N__36599\
        );

    \I__7604\ : InMux
    port map (
            O => \N__36604\,
            I => \N__36596\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__36599\,
            I => \N__36593\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__36596\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__36593\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__7600\ : CascadeMux
    port map (
            O => \N__36588\,
            I => \N__36585\
        );

    \I__7599\ : InMux
    port map (
            O => \N__36585\,
            I => \N__36582\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__36582\,
            I => \N__36579\
        );

    \I__7597\ : Span4Mux_v
    port map (
            O => \N__36579\,
            I => \N__36576\
        );

    \I__7596\ : Odrv4
    port map (
            O => \N__36576\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__7595\ : CascadeMux
    port map (
            O => \N__36573\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\
        );

    \I__7594\ : InMux
    port map (
            O => \N__36570\,
            I => \N__36564\
        );

    \I__7593\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36564\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__36564\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__36561\,
            I => \N__36558\
        );

    \I__7590\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36552\
        );

    \I__7589\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36552\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__36552\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__7587\ : InMux
    port map (
            O => \N__36549\,
            I => \N__36546\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__36546\,
            I => \N__36543\
        );

    \I__7585\ : Odrv4
    port map (
            O => \N__36543\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__7584\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36536\
        );

    \I__7583\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36532\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__36536\,
            I => \N__36529\
        );

    \I__7581\ : InMux
    port map (
            O => \N__36535\,
            I => \N__36526\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__36532\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__7579\ : Odrv4
    port map (
            O => \N__36529\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__36526\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__7577\ : InMux
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__36516\,
            I => \N__36510\
        );

    \I__7575\ : InMux
    port map (
            O => \N__36515\,
            I => \N__36507\
        );

    \I__7574\ : InMux
    port map (
            O => \N__36514\,
            I => \N__36502\
        );

    \I__7573\ : InMux
    port map (
            O => \N__36513\,
            I => \N__36502\
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__36510\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__36507\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__36502\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__7569\ : InMux
    port map (
            O => \N__36495\,
            I => \N__36492\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__36492\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__7567\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36485\
        );

    \I__7566\ : InMux
    port map (
            O => \N__36488\,
            I => \N__36481\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__36485\,
            I => \N__36478\
        );

    \I__7564\ : InMux
    port map (
            O => \N__36484\,
            I => \N__36475\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__36481\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__7562\ : Odrv4
    port map (
            O => \N__36478\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__36475\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__7560\ : InMux
    port map (
            O => \N__36468\,
            I => \N__36464\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36461\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36464\,
            I => \N__36454\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__36461\,
            I => \N__36454\
        );

    \I__7556\ : InMux
    port map (
            O => \N__36460\,
            I => \N__36451\
        );

    \I__7555\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36448\
        );

    \I__7554\ : Span4Mux_v
    port map (
            O => \N__36454\,
            I => \N__36441\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N__36441\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36448\,
            I => \N__36441\
        );

    \I__7551\ : Odrv4
    port map (
            O => \N__36441\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__7550\ : CascadeMux
    port map (
            O => \N__36438\,
            I => \N__36435\
        );

    \I__7549\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__36432\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__7547\ : InMux
    port map (
            O => \N__36429\,
            I => \N__36425\
        );

    \I__7546\ : InMux
    port map (
            O => \N__36428\,
            I => \N__36421\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36425\,
            I => \N__36418\
        );

    \I__7544\ : InMux
    port map (
            O => \N__36424\,
            I => \N__36415\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__36421\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__7542\ : Odrv4
    port map (
            O => \N__36418\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__36415\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__7540\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36404\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36401\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__36404\,
            I => \N__36394\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__36401\,
            I => \N__36394\
        );

    \I__7536\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36389\
        );

    \I__7535\ : InMux
    port map (
            O => \N__36399\,
            I => \N__36389\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__36394\,
            I => \N__36384\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__36389\,
            I => \N__36384\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__36384\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__7531\ : InMux
    port map (
            O => \N__36381\,
            I => \N__36378\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__36378\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__36375\,
            I => \N__36372\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36372\,
            I => \N__36366\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36371\,
            I => \N__36363\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36370\,
            I => \N__36358\
        );

    \I__7525\ : InMux
    port map (
            O => \N__36369\,
            I => \N__36358\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__36366\,
            I => \N__36355\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__36363\,
            I => \N__36352\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__36358\,
            I => \N__36349\
        );

    \I__7521\ : Span4Mux_h
    port map (
            O => \N__36355\,
            I => \N__36346\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__36352\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__7519\ : Odrv4
    port map (
            O => \N__36349\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__7518\ : Odrv4
    port map (
            O => \N__36346\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__7517\ : InMux
    port map (
            O => \N__36339\,
            I => \N__36336\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__36336\,
            I => \N__36333\
        );

    \I__7515\ : Span4Mux_h
    port map (
            O => \N__36333\,
            I => \N__36329\
        );

    \I__7514\ : InMux
    port map (
            O => \N__36332\,
            I => \N__36326\
        );

    \I__7513\ : Odrv4
    port map (
            O => \N__36329\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__36326\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__7511\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36315\
        );

    \I__7510\ : InMux
    port map (
            O => \N__36320\,
            I => \N__36315\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__36315\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__7508\ : InMux
    port map (
            O => \N__36312\,
            I => \N__36309\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__36306\,
            I => \N__36302\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36305\,
            I => \N__36299\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__36302\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__36299\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__7502\ : InMux
    port map (
            O => \N__36294\,
            I => \N__36289\
        );

    \I__7501\ : InMux
    port map (
            O => \N__36293\,
            I => \N__36284\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36292\,
            I => \N__36284\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__36289\,
            I => \N__36280\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36284\,
            I => \N__36277\
        );

    \I__7497\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36274\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__36280\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__36277\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__36274\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__7493\ : CascadeMux
    port map (
            O => \N__36267\,
            I => \N__36264\
        );

    \I__7492\ : InMux
    port map (
            O => \N__36264\,
            I => \N__36258\
        );

    \I__7491\ : InMux
    port map (
            O => \N__36263\,
            I => \N__36258\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__36258\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__7489\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36251\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36248\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__36251\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__36248\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__7485\ : InMux
    port map (
            O => \N__36243\,
            I => \N__36240\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36240\,
            I => \N__36237\
        );

    \I__7483\ : Span4Mux_v
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__7482\ : Odrv4
    port map (
            O => \N__36234\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__36231\,
            I => \N__36227\
        );

    \I__7480\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36224\
        );

    \I__7479\ : InMux
    port map (
            O => \N__36227\,
            I => \N__36221\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__36224\,
            I => \N__36217\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36221\,
            I => \N__36214\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36211\
        );

    \I__7475\ : Odrv4
    port map (
            O => \N__36217\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__36214\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7473\ : LocalMux
    port map (
            O => \N__36211\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__7472\ : CEMux
    port map (
            O => \N__36204\,
            I => \N__36200\
        );

    \I__7471\ : CEMux
    port map (
            O => \N__36203\,
            I => \N__36197\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__36200\,
            I => \N__36191\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__36197\,
            I => \N__36188\
        );

    \I__7468\ : CEMux
    port map (
            O => \N__36196\,
            I => \N__36185\
        );

    \I__7467\ : CEMux
    port map (
            O => \N__36195\,
            I => \N__36182\
        );

    \I__7466\ : CEMux
    port map (
            O => \N__36194\,
            I => \N__36179\
        );

    \I__7465\ : Span4Mux_v
    port map (
            O => \N__36191\,
            I => \N__36175\
        );

    \I__7464\ : Span4Mux_h
    port map (
            O => \N__36188\,
            I => \N__36172\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__36185\,
            I => \N__36169\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__36182\,
            I => \N__36166\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__36179\,
            I => \N__36163\
        );

    \I__7460\ : CEMux
    port map (
            O => \N__36178\,
            I => \N__36160\
        );

    \I__7459\ : Span4Mux_v
    port map (
            O => \N__36175\,
            I => \N__36157\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__36172\,
            I => \N__36154\
        );

    \I__7457\ : Span4Mux_v
    port map (
            O => \N__36169\,
            I => \N__36145\
        );

    \I__7456\ : Span4Mux_v
    port map (
            O => \N__36166\,
            I => \N__36145\
        );

    \I__7455\ : Span4Mux_h
    port map (
            O => \N__36163\,
            I => \N__36145\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36160\,
            I => \N__36145\
        );

    \I__7453\ : Span4Mux_v
    port map (
            O => \N__36157\,
            I => \N__36142\
        );

    \I__7452\ : Span4Mux_v
    port map (
            O => \N__36154\,
            I => \N__36139\
        );

    \I__7451\ : Span4Mux_v
    port map (
            O => \N__36145\,
            I => \N__36136\
        );

    \I__7450\ : Span4Mux_v
    port map (
            O => \N__36142\,
            I => \N__36133\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__36139\,
            I => \N__36130\
        );

    \I__7448\ : Span4Mux_v
    port map (
            O => \N__36136\,
            I => \N__36127\
        );

    \I__7447\ : Odrv4
    port map (
            O => \N__36133\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7446\ : Odrv4
    port map (
            O => \N__36130\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__36127\,
            I => \delay_measurement_inst.delay_tr_timer.N_200_i\
        );

    \I__7444\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36114\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36119\,
            I => \N__36114\
        );

    \I__7442\ : LocalMux
    port map (
            O => \N__36114\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__7441\ : CascadeMux
    port map (
            O => \N__36111\,
            I => \N__36108\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36102\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36107\,
            I => \N__36102\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__36102\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36099\,
            I => \N__36096\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__36093\
        );

    \I__7435\ : Odrv4
    port map (
            O => \N__36093\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__7434\ : CascadeMux
    port map (
            O => \N__36090\,
            I => \N__36085\
        );

    \I__7433\ : InMux
    port map (
            O => \N__36089\,
            I => \N__36082\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36070\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36070\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36082\,
            I => \N__36067\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36081\,
            I => \N__36052\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36080\,
            I => \N__36052\
        );

    \I__7427\ : InMux
    port map (
            O => \N__36079\,
            I => \N__36052\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36052\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36077\,
            I => \N__36052\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36052\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36075\,
            I => \N__36052\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__36070\,
            I => \N__36049\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__36067\,
            I => \N__36044\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__36052\,
            I => \N__36044\
        );

    \I__7419\ : Span4Mux_h
    port map (
            O => \N__36049\,
            I => \N__36041\
        );

    \I__7418\ : Span4Mux_h
    port map (
            O => \N__36044\,
            I => \N__36038\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__36041\,
            I => \N__36035\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__36038\,
            I => \N__36032\
        );

    \I__7415\ : Span4Mux_h
    port map (
            O => \N__36035\,
            I => \N__36029\
        );

    \I__7414\ : Span4Mux_h
    port map (
            O => \N__36032\,
            I => \N__36026\
        );

    \I__7413\ : Odrv4
    port map (
            O => \N__36029\,
            I => \pwm_generator_inst.N_16\
        );

    \I__7412\ : Odrv4
    port map (
            O => \N__36026\,
            I => \pwm_generator_inst.N_16\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36021\,
            I => \N__35993\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36020\,
            I => \N__35993\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36019\,
            I => \N__35986\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36018\,
            I => \N__35986\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36017\,
            I => \N__35986\
        );

    \I__7406\ : InMux
    port map (
            O => \N__36016\,
            I => \N__35969\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36015\,
            I => \N__35969\
        );

    \I__7404\ : InMux
    port map (
            O => \N__36014\,
            I => \N__35969\
        );

    \I__7403\ : InMux
    port map (
            O => \N__36013\,
            I => \N__35969\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36012\,
            I => \N__35969\
        );

    \I__7401\ : InMux
    port map (
            O => \N__36011\,
            I => \N__35969\
        );

    \I__7400\ : InMux
    port map (
            O => \N__36010\,
            I => \N__35969\
        );

    \I__7399\ : InMux
    port map (
            O => \N__36009\,
            I => \N__35969\
        );

    \I__7398\ : InMux
    port map (
            O => \N__36008\,
            I => \N__35954\
        );

    \I__7397\ : InMux
    port map (
            O => \N__36007\,
            I => \N__35954\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36006\,
            I => \N__35954\
        );

    \I__7395\ : InMux
    port map (
            O => \N__36005\,
            I => \N__35954\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36004\,
            I => \N__35954\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36003\,
            I => \N__35954\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36002\,
            I => \N__35954\
        );

    \I__7391\ : CascadeMux
    port map (
            O => \N__36001\,
            I => \N__35947\
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__36000\,
            I => \N__35944\
        );

    \I__7389\ : CascadeMux
    port map (
            O => \N__35999\,
            I => \N__35940\
        );

    \I__7388\ : CascadeMux
    port map (
            O => \N__35998\,
            I => \N__35936\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__35993\,
            I => \N__35931\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__35986\,
            I => \N__35931\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__35969\,
            I => \N__35926\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__35954\,
            I => \N__35926\
        );

    \I__7383\ : InMux
    port map (
            O => \N__35953\,
            I => \N__35921\
        );

    \I__7382\ : InMux
    port map (
            O => \N__35952\,
            I => \N__35921\
        );

    \I__7381\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35906\
        );

    \I__7380\ : InMux
    port map (
            O => \N__35950\,
            I => \N__35906\
        );

    \I__7379\ : InMux
    port map (
            O => \N__35947\,
            I => \N__35906\
        );

    \I__7378\ : InMux
    port map (
            O => \N__35944\,
            I => \N__35906\
        );

    \I__7377\ : InMux
    port map (
            O => \N__35943\,
            I => \N__35906\
        );

    \I__7376\ : InMux
    port map (
            O => \N__35940\,
            I => \N__35906\
        );

    \I__7375\ : InMux
    port map (
            O => \N__35939\,
            I => \N__35906\
        );

    \I__7374\ : InMux
    port map (
            O => \N__35936\,
            I => \N__35903\
        );

    \I__7373\ : Span4Mux_v
    port map (
            O => \N__35931\,
            I => \N__35899\
        );

    \I__7372\ : Span4Mux_v
    port map (
            O => \N__35926\,
            I => \N__35896\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__35921\,
            I => \N__35893\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__35906\,
            I => \N__35888\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__35903\,
            I => \N__35888\
        );

    \I__7368\ : CascadeMux
    port map (
            O => \N__35902\,
            I => \N__35885\
        );

    \I__7367\ : Span4Mux_h
    port map (
            O => \N__35899\,
            I => \N__35881\
        );

    \I__7366\ : Sp12to4
    port map (
            O => \N__35896\,
            I => \N__35878\
        );

    \I__7365\ : Span4Mux_h
    port map (
            O => \N__35893\,
            I => \N__35875\
        );

    \I__7364\ : Span4Mux_h
    port map (
            O => \N__35888\,
            I => \N__35872\
        );

    \I__7363\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35867\
        );

    \I__7362\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35867\
        );

    \I__7361\ : Sp12to4
    port map (
            O => \N__35881\,
            I => \N__35862\
        );

    \I__7360\ : Span12Mux_s8_h
    port map (
            O => \N__35878\,
            I => \N__35862\
        );

    \I__7359\ : Odrv4
    port map (
            O => \N__35875\,
            I => \N_19_1\
        );

    \I__7358\ : Odrv4
    port map (
            O => \N__35872\,
            I => \N_19_1\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__35867\,
            I => \N_19_1\
        );

    \I__7356\ : Odrv12
    port map (
            O => \N__35862\,
            I => \N_19_1\
        );

    \I__7355\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35847\
        );

    \I__7354\ : InMux
    port map (
            O => \N__35852\,
            I => \N__35847\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35843\
        );

    \I__7352\ : InMux
    port map (
            O => \N__35846\,
            I => \N__35833\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__35843\,
            I => \N__35830\
        );

    \I__7350\ : InMux
    port map (
            O => \N__35842\,
            I => \N__35815\
        );

    \I__7349\ : InMux
    port map (
            O => \N__35841\,
            I => \N__35815\
        );

    \I__7348\ : InMux
    port map (
            O => \N__35840\,
            I => \N__35815\
        );

    \I__7347\ : InMux
    port map (
            O => \N__35839\,
            I => \N__35815\
        );

    \I__7346\ : InMux
    port map (
            O => \N__35838\,
            I => \N__35815\
        );

    \I__7345\ : InMux
    port map (
            O => \N__35837\,
            I => \N__35815\
        );

    \I__7344\ : InMux
    port map (
            O => \N__35836\,
            I => \N__35815\
        );

    \I__7343\ : LocalMux
    port map (
            O => \N__35833\,
            I => \N__35812\
        );

    \I__7342\ : Sp12to4
    port map (
            O => \N__35830\,
            I => \N__35805\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__35815\,
            I => \N__35805\
        );

    \I__7340\ : Sp12to4
    port map (
            O => \N__35812\,
            I => \N__35805\
        );

    \I__7339\ : Odrv12
    port map (
            O => \N__35805\,
            I => \pwm_generator_inst.N_17\
        );

    \I__7338\ : CascadeMux
    port map (
            O => \N__35802\,
            I => \N__35799\
        );

    \I__7337\ : InMux
    port map (
            O => \N__35799\,
            I => \N__35796\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35793\
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__35793\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__7334\ : InMux
    port map (
            O => \N__35790\,
            I => \N__35787\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__35787\,
            I => \N__35783\
        );

    \I__7332\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35780\
        );

    \I__7331\ : Span12Mux_h
    port map (
            O => \N__35783\,
            I => \N__35777\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__35780\,
            I => \N__35774\
        );

    \I__7329\ : Odrv12
    port map (
            O => \N__35777\,
            I => state_ns_i_a3_1
        );

    \I__7328\ : Odrv4
    port map (
            O => \N__35774\,
            I => state_ns_i_a3_1
        );

    \I__7327\ : IoInMux
    port map (
            O => \N__35769\,
            I => \N__35766\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__35766\,
            I => \N__35763\
        );

    \I__7325\ : IoSpan4Mux
    port map (
            O => \N__35763\,
            I => \N__35760\
        );

    \I__7324\ : Span4Mux_s1_v
    port map (
            O => \N__35760\,
            I => \N__35757\
        );

    \I__7323\ : Sp12to4
    port map (
            O => \N__35757\,
            I => \N__35754\
        );

    \I__7322\ : Span12Mux_v
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__7321\ : Span12Mux_v
    port map (
            O => \N__35751\,
            I => \N__35747\
        );

    \I__7320\ : InMux
    port map (
            O => \N__35750\,
            I => \N__35744\
        );

    \I__7319\ : Odrv12
    port map (
            O => \N__35747\,
            I => \T45_c\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__35744\,
            I => \T45_c\
        );

    \I__7317\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35735\
        );

    \I__7316\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35732\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__35735\,
            I => \N__35726\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__35732\,
            I => \N__35726\
        );

    \I__7313\ : InMux
    port map (
            O => \N__35731\,
            I => \N__35723\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__35726\,
            I => \N__35718\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__35723\,
            I => \N__35718\
        );

    \I__7310\ : Span4Mux_h
    port map (
            O => \N__35718\,
            I => \N__35715\
        );

    \I__7309\ : Span4Mux_h
    port map (
            O => \N__35715\,
            I => \N__35712\
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__35712\,
            I => il_min_comp2_c
        );

    \I__7307\ : InMux
    port map (
            O => \N__35709\,
            I => \N__35705\
        );

    \I__7306\ : InMux
    port map (
            O => \N__35708\,
            I => \N__35702\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__35705\,
            I => \N__35699\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__35702\,
            I => \N__35696\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__35699\,
            I => \N__35691\
        );

    \I__7302\ : Span4Mux_v
    port map (
            O => \N__35696\,
            I => \N__35691\
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__35691\,
            I => \phase_controller_inst2.time_passed_RNIG7JF\
        );

    \I__7300\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35685\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__35685\,
            I => \N__35682\
        );

    \I__7298\ : Span4Mux_v
    port map (
            O => \N__35682\,
            I => \N__35679\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__35679\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__7296\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35672\
        );

    \I__7295\ : InMux
    port map (
            O => \N__35675\,
            I => \N__35665\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__35672\,
            I => \N__35654\
        );

    \I__7293\ : InMux
    port map (
            O => \N__35671\,
            I => \N__35651\
        );

    \I__7292\ : InMux
    port map (
            O => \N__35670\,
            I => \N__35646\
        );

    \I__7291\ : InMux
    port map (
            O => \N__35669\,
            I => \N__35646\
        );

    \I__7290\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35643\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35637\
        );

    \I__7288\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35634\
        );

    \I__7287\ : InMux
    port map (
            O => \N__35663\,
            I => \N__35627\
        );

    \I__7286\ : InMux
    port map (
            O => \N__35662\,
            I => \N__35627\
        );

    \I__7285\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35627\
        );

    \I__7284\ : InMux
    port map (
            O => \N__35660\,
            I => \N__35618\
        );

    \I__7283\ : InMux
    port map (
            O => \N__35659\,
            I => \N__35618\
        );

    \I__7282\ : InMux
    port map (
            O => \N__35658\,
            I => \N__35618\
        );

    \I__7281\ : InMux
    port map (
            O => \N__35657\,
            I => \N__35618\
        );

    \I__7280\ : Span4Mux_v
    port map (
            O => \N__35654\,
            I => \N__35611\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__35651\,
            I => \N__35611\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__35646\,
            I => \N__35611\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__35643\,
            I => \N__35608\
        );

    \I__7276\ : InMux
    port map (
            O => \N__35642\,
            I => \N__35604\
        );

    \I__7275\ : InMux
    port map (
            O => \N__35641\,
            I => \N__35601\
        );

    \I__7274\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35598\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__35637\,
            I => \N__35572\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__35634\,
            I => \N__35572\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__35627\,
            I => \N__35572\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__35618\,
            I => \N__35572\
        );

    \I__7269\ : Span4Mux_v
    port map (
            O => \N__35611\,
            I => \N__35569\
        );

    \I__7268\ : Span4Mux_v
    port map (
            O => \N__35608\,
            I => \N__35566\
        );

    \I__7267\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35563\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35560\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__35601\,
            I => \N__35555\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__35598\,
            I => \N__35555\
        );

    \I__7263\ : InMux
    port map (
            O => \N__35597\,
            I => \N__35548\
        );

    \I__7262\ : InMux
    port map (
            O => \N__35596\,
            I => \N__35548\
        );

    \I__7261\ : InMux
    port map (
            O => \N__35595\,
            I => \N__35548\
        );

    \I__7260\ : InMux
    port map (
            O => \N__35594\,
            I => \N__35539\
        );

    \I__7259\ : InMux
    port map (
            O => \N__35593\,
            I => \N__35539\
        );

    \I__7258\ : InMux
    port map (
            O => \N__35592\,
            I => \N__35539\
        );

    \I__7257\ : InMux
    port map (
            O => \N__35591\,
            I => \N__35539\
        );

    \I__7256\ : CascadeMux
    port map (
            O => \N__35590\,
            I => \N__35534\
        );

    \I__7255\ : CascadeMux
    port map (
            O => \N__35589\,
            I => \N__35530\
        );

    \I__7254\ : CascadeMux
    port map (
            O => \N__35588\,
            I => \N__35526\
        );

    \I__7253\ : CascadeMux
    port map (
            O => \N__35587\,
            I => \N__35521\
        );

    \I__7252\ : CascadeMux
    port map (
            O => \N__35586\,
            I => \N__35517\
        );

    \I__7251\ : CascadeMux
    port map (
            O => \N__35585\,
            I => \N__35513\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__35584\,
            I => \N__35509\
        );

    \I__7249\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35495\
        );

    \I__7248\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35495\
        );

    \I__7247\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35492\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__35572\,
            I => \N__35489\
        );

    \I__7245\ : Span4Mux_v
    port map (
            O => \N__35569\,
            I => \N__35484\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__35566\,
            I => \N__35484\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__35563\,
            I => \N__35481\
        );

    \I__7242\ : Span4Mux_v
    port map (
            O => \N__35560\,
            I => \N__35472\
        );

    \I__7241\ : Span4Mux_v
    port map (
            O => \N__35555\,
            I => \N__35472\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35472\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__35539\,
            I => \N__35472\
        );

    \I__7238\ : CascadeMux
    port map (
            O => \N__35538\,
            I => \N__35468\
        );

    \I__7237\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35452\
        );

    \I__7236\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35452\
        );

    \I__7235\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35452\
        );

    \I__7234\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35452\
        );

    \I__7233\ : InMux
    port map (
            O => \N__35529\,
            I => \N__35452\
        );

    \I__7232\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35452\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35525\,
            I => \N__35452\
        );

    \I__7230\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35435\
        );

    \I__7229\ : InMux
    port map (
            O => \N__35521\,
            I => \N__35435\
        );

    \I__7228\ : InMux
    port map (
            O => \N__35520\,
            I => \N__35435\
        );

    \I__7227\ : InMux
    port map (
            O => \N__35517\,
            I => \N__35435\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35435\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35435\
        );

    \I__7224\ : InMux
    port map (
            O => \N__35512\,
            I => \N__35435\
        );

    \I__7223\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35435\
        );

    \I__7222\ : InMux
    port map (
            O => \N__35508\,
            I => \N__35430\
        );

    \I__7221\ : InMux
    port map (
            O => \N__35507\,
            I => \N__35430\
        );

    \I__7220\ : CascadeMux
    port map (
            O => \N__35506\,
            I => \N__35427\
        );

    \I__7219\ : CascadeMux
    port map (
            O => \N__35505\,
            I => \N__35423\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__35504\,
            I => \N__35419\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__35503\,
            I => \N__35415\
        );

    \I__7216\ : CascadeMux
    port map (
            O => \N__35502\,
            I => \N__35410\
        );

    \I__7215\ : CascadeMux
    port map (
            O => \N__35501\,
            I => \N__35406\
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__35500\,
            I => \N__35402\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35495\,
            I => \N__35396\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__35492\,
            I => \N__35396\
        );

    \I__7211\ : Span4Mux_h
    port map (
            O => \N__35489\,
            I => \N__35393\
        );

    \I__7210\ : Span4Mux_v
    port map (
            O => \N__35484\,
            I => \N__35386\
        );

    \I__7209\ : Span4Mux_v
    port map (
            O => \N__35481\,
            I => \N__35386\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__35472\,
            I => \N__35386\
        );

    \I__7207\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35379\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35379\
        );

    \I__7205\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35379\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__35452\,
            I => \N__35372\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__35435\,
            I => \N__35372\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__35430\,
            I => \N__35372\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35427\,
            I => \N__35355\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35355\
        );

    \I__7199\ : InMux
    port map (
            O => \N__35423\,
            I => \N__35355\
        );

    \I__7198\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35355\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35419\,
            I => \N__35355\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35418\,
            I => \N__35355\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35415\,
            I => \N__35355\
        );

    \I__7194\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35355\
        );

    \I__7193\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35340\
        );

    \I__7192\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35340\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35340\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35406\,
            I => \N__35340\
        );

    \I__7189\ : InMux
    port map (
            O => \N__35405\,
            I => \N__35340\
        );

    \I__7188\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35340\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35340\
        );

    \I__7186\ : Span12Mux_s11_h
    port map (
            O => \N__35396\,
            I => \N__35337\
        );

    \I__7185\ : Span4Mux_h
    port map (
            O => \N__35393\,
            I => \N__35334\
        );

    \I__7184\ : Span4Mux_h
    port map (
            O => \N__35386\,
            I => \N__35331\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__35379\,
            I => \N__35328\
        );

    \I__7182\ : Span4Mux_v
    port map (
            O => \N__35372\,
            I => \N__35321\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__35355\,
            I => \N__35321\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35340\,
            I => \N__35321\
        );

    \I__7179\ : Span12Mux_v
    port map (
            O => \N__35337\,
            I => \N__35318\
        );

    \I__7178\ : Span4Mux_h
    port map (
            O => \N__35334\,
            I => \N__35313\
        );

    \I__7177\ : Span4Mux_h
    port map (
            O => \N__35331\,
            I => \N__35313\
        );

    \I__7176\ : Span4Mux_v
    port map (
            O => \N__35328\,
            I => \N__35308\
        );

    \I__7175\ : Span4Mux_v
    port map (
            O => \N__35321\,
            I => \N__35308\
        );

    \I__7174\ : Odrv12
    port map (
            O => \N__35318\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7173\ : Odrv4
    port map (
            O => \N__35313\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7172\ : Odrv4
    port map (
            O => \N__35308\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7171\ : InMux
    port map (
            O => \N__35301\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__7170\ : InMux
    port map (
            O => \N__35298\,
            I => \N__35291\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35291\
        );

    \I__7168\ : CascadeMux
    port map (
            O => \N__35296\,
            I => \N__35279\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__35291\,
            I => \N__35273\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35258\
        );

    \I__7165\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35258\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35258\
        );

    \I__7163\ : InMux
    port map (
            O => \N__35287\,
            I => \N__35258\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35286\,
            I => \N__35258\
        );

    \I__7161\ : InMux
    port map (
            O => \N__35285\,
            I => \N__35258\
        );

    \I__7160\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35258\
        );

    \I__7159\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35253\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35282\,
            I => \N__35253\
        );

    \I__7157\ : InMux
    port map (
            O => \N__35279\,
            I => \N__35250\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35278\,
            I => \N__35243\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35243\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35243\
        );

    \I__7153\ : Span4Mux_h
    port map (
            O => \N__35273\,
            I => \N__35238\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35258\,
            I => \N__35238\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__35253\,
            I => \N__35235\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35250\,
            I => \N__35230\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__35243\,
            I => \N__35230\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__35238\,
            I => \N__35227\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__35235\,
            I => \N__35224\
        );

    \I__7146\ : Span4Mux_h
    port map (
            O => \N__35230\,
            I => \N__35219\
        );

    \I__7145\ : Span4Mux_v
    port map (
            O => \N__35227\,
            I => \N__35219\
        );

    \I__7144\ : Odrv4
    port map (
            O => \N__35224\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__35219\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__7142\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__35211\,
            I => \N__35205\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35202\
        );

    \I__7139\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35197\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35197\
        );

    \I__7137\ : Span12Mux_v
    port map (
            O => \N__35205\,
            I => \N__35194\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__35202\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__35197\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7134\ : Odrv12
    port map (
            O => \N__35194\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__7133\ : InMux
    port map (
            O => \N__35187\,
            I => \N__35183\
        );

    \I__7132\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35179\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__35183\,
            I => \N__35176\
        );

    \I__7130\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35173\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35179\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__7128\ : Odrv4
    port map (
            O => \N__35176\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35173\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__7126\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35162\
        );

    \I__7125\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35158\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__35162\,
            I => \N__35155\
        );

    \I__7123\ : InMux
    port map (
            O => \N__35161\,
            I => \N__35152\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35158\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__35155\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35152\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__7119\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35140\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35137\
        );

    \I__7117\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35134\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35131\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__35137\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35134\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__7113\ : Odrv4
    port map (
            O => \N__35131\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__7112\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35120\
        );

    \I__7111\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35116\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__35120\,
            I => \N__35113\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35110\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__35116\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__35113\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__7106\ : LocalMux
    port map (
            O => \N__35110\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35103\,
            I => \N__35099\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35102\,
            I => \N__35095\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__35099\,
            I => \N__35092\
        );

    \I__7102\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35089\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__35095\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__7100\ : Odrv4
    port map (
            O => \N__35092\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__35089\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35077\
        );

    \I__7097\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35074\
        );

    \I__7096\ : InMux
    port map (
            O => \N__35080\,
            I => \N__35071\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35077\,
            I => \N__35068\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__35074\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35071\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__7092\ : Odrv4
    port map (
            O => \N__35068\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__7091\ : InMux
    port map (
            O => \N__35061\,
            I => \N__35056\
        );

    \I__7090\ : InMux
    port map (
            O => \N__35060\,
            I => \N__35053\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35059\,
            I => \N__35050\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__35056\,
            I => \N__35047\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__35053\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35050\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__7085\ : Odrv4
    port map (
            O => \N__35047\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__7084\ : CascadeMux
    port map (
            O => \N__35040\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35032\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35029\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35026\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__35032\,
            I => \N__35023\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__35029\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__35026\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__35023\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35016\,
            I => \N__35013\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__35013\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35010\,
            I => \N__35005\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35009\,
            I => \N__35002\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35008\,
            I => \N__34999\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__35005\,
            I => \N__34996\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35002\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__34999\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__7068\ : Odrv4
    port map (
            O => \N__34996\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__7067\ : CascadeMux
    port map (
            O => \N__34989\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__7066\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34981\
        );

    \I__7065\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34978\
        );

    \I__7064\ : InMux
    port map (
            O => \N__34984\,
            I => \N__34975\
        );

    \I__7063\ : LocalMux
    port map (
            O => \N__34981\,
            I => \N__34972\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__34978\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__34975\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__34972\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__7059\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34947\
        );

    \I__7058\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34947\
        );

    \I__7057\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34947\
        );

    \I__7056\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34947\
        );

    \I__7055\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34942\
        );

    \I__7054\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34942\
        );

    \I__7053\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34933\
        );

    \I__7052\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34933\
        );

    \I__7051\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34933\
        );

    \I__7050\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34933\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__34947\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__34942\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__34933\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__7046\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__7045\ : LocalMux
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__7044\ : Odrv4
    port map (
            O => \N__34920\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__7043\ : InMux
    port map (
            O => \N__34917\,
            I => \N__34914\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__34914\,
            I => \N__34911\
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__34911\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__7040\ : CascadeMux
    port map (
            O => \N__34908\,
            I => \N__34905\
        );

    \I__7039\ : InMux
    port map (
            O => \N__34905\,
            I => \N__34902\
        );

    \I__7038\ : LocalMux
    port map (
            O => \N__34902\,
            I => \N__34899\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__34899\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__7036\ : CascadeMux
    port map (
            O => \N__34896\,
            I => \N__34893\
        );

    \I__7035\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34890\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__34890\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__7033\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34884\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__34884\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__7031\ : InMux
    port map (
            O => \N__34881\,
            I => \N__34878\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__34878\,
            I => \N__34875\
        );

    \I__7029\ : Odrv4
    port map (
            O => \N__34875\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__7028\ : CascadeMux
    port map (
            O => \N__34872\,
            I => \N__34869\
        );

    \I__7027\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34866\
        );

    \I__7026\ : LocalMux
    port map (
            O => \N__34866\,
            I => \N__34863\
        );

    \I__7025\ : Odrv4
    port map (
            O => \N__34863\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__7024\ : CascadeMux
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__7023\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34854\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__34854\,
            I => \N__34851\
        );

    \I__7021\ : Odrv4
    port map (
            O => \N__34851\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__7020\ : InMux
    port map (
            O => \N__34848\,
            I => \N__34845\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__34845\,
            I => \N__34842\
        );

    \I__7018\ : Odrv12
    port map (
            O => \N__34842\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__7017\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34836\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__34836\,
            I => \N__34833\
        );

    \I__7015\ : Span4Mux_h
    port map (
            O => \N__34833\,
            I => \N__34830\
        );

    \I__7014\ : Odrv4
    port map (
            O => \N__34830\,
            I => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\
        );

    \I__7013\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34824\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__34824\,
            I => \N__34821\
        );

    \I__7011\ : Span4Mux_h
    port map (
            O => \N__34821\,
            I => \N__34818\
        );

    \I__7010\ : Odrv4
    port map (
            O => \N__34818\,
            I => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\
        );

    \I__7009\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34812\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__34812\,
            I => \N__34809\
        );

    \I__7007\ : Span4Mux_v
    port map (
            O => \N__34809\,
            I => \N__34806\
        );

    \I__7006\ : Odrv4
    port map (
            O => \N__34806\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__7005\ : InMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__34800\,
            I => \N__34797\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__34797\,
            I => \N__34794\
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__34794\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__7001\ : CascadeMux
    port map (
            O => \N__34791\,
            I => \N__34788\
        );

    \I__7000\ : InMux
    port map (
            O => \N__34788\,
            I => \N__34785\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__34785\,
            I => \N__34782\
        );

    \I__6998\ : Span4Mux_h
    port map (
            O => \N__34782\,
            I => \N__34779\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__34779\,
            I => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\
        );

    \I__6996\ : CascadeMux
    port map (
            O => \N__34776\,
            I => \N__34773\
        );

    \I__6995\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34770\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__34770\,
            I => \N__34767\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__34767\,
            I => \N__34764\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__34764\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__34761\,
            I => \N__34758\
        );

    \I__6990\ : InMux
    port map (
            O => \N__34758\,
            I => \N__34754\
        );

    \I__6989\ : InMux
    port map (
            O => \N__34757\,
            I => \N__34751\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__34754\,
            I => \N__34748\
        );

    \I__6987\ : LocalMux
    port map (
            O => \N__34751\,
            I => \N__34745\
        );

    \I__6986\ : Span4Mux_v
    port map (
            O => \N__34748\,
            I => \N__34742\
        );

    \I__6985\ : Odrv12
    port map (
            O => \N__34745\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__34742\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__6983\ : InMux
    port map (
            O => \N__34737\,
            I => \N__34734\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__6981\ : Odrv12
    port map (
            O => \N__34731\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__6980\ : CascadeMux
    port map (
            O => \N__34728\,
            I => \N__34725\
        );

    \I__6979\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34722\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__34722\,
            I => \N__34719\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__34719\,
            I => \N__34716\
        );

    \I__6976\ : Odrv4
    port map (
            O => \N__34716\,
            I => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__34713\,
            I => \N__34710\
        );

    \I__6974\ : InMux
    port map (
            O => \N__34710\,
            I => \N__34707\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__34707\,
            I => \N__34704\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__34704\,
            I => \N__34701\
        );

    \I__6971\ : Odrv4
    port map (
            O => \N__34701\,
            I => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\
        );

    \I__6970\ : InMux
    port map (
            O => \N__34698\,
            I => \N__34695\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__34695\,
            I => \N__34692\
        );

    \I__6968\ : Span4Mux_v
    port map (
            O => \N__34692\,
            I => \N__34689\
        );

    \I__6967\ : Odrv4
    port map (
            O => \N__34689\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__34686\,
            I => \N__34683\
        );

    \I__6965\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34680\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__34677\,
            I => \N__34674\
        );

    \I__6962\ : Odrv4
    port map (
            O => \N__34674\,
            I => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\
        );

    \I__6961\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34668\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__34668\,
            I => \N__34665\
        );

    \I__6959\ : Span4Mux_v
    port map (
            O => \N__34665\,
            I => \N__34662\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__34662\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__6957\ : CascadeMux
    port map (
            O => \N__34659\,
            I => \N__34656\
        );

    \I__6956\ : InMux
    port map (
            O => \N__34656\,
            I => \N__34653\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__34653\,
            I => \N__34650\
        );

    \I__6954\ : Span4Mux_v
    port map (
            O => \N__34650\,
            I => \N__34647\
        );

    \I__6953\ : Odrv4
    port map (
            O => \N__34647\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__6952\ : InMux
    port map (
            O => \N__34644\,
            I => \N__34641\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__34641\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\
        );

    \I__6950\ : InMux
    port map (
            O => \N__34638\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_28\
        );

    \I__6949\ : InMux
    port map (
            O => \N__34635\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__6948\ : CascadeMux
    port map (
            O => \N__34632\,
            I => \N__34629\
        );

    \I__6947\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34626\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__34626\,
            I => \N__34623\
        );

    \I__6945\ : Span4Mux_v
    port map (
            O => \N__34623\,
            I => \N__34620\
        );

    \I__6944\ : Odrv4
    port map (
            O => \N__34620\,
            I => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\
        );

    \I__6943\ : CascadeMux
    port map (
            O => \N__34617\,
            I => \N__34614\
        );

    \I__6942\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34611\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__34611\,
            I => \N__34608\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__34608\,
            I => \N__34605\
        );

    \I__6939\ : Odrv4
    port map (
            O => \N__34605\,
            I => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__34602\,
            I => \N__34599\
        );

    \I__6937\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34596\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__34596\,
            I => \N__34593\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__34593\,
            I => \N__34590\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__34590\,
            I => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\
        );

    \I__6933\ : CascadeMux
    port map (
            O => \N__34587\,
            I => \N__34584\
        );

    \I__6932\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34581\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__34581\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__6930\ : CascadeMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__6929\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34572\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__34572\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__6927\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34566\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__34566\,
            I => \N__34563\
        );

    \I__6925\ : Odrv4
    port map (
            O => \N__34563\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__6924\ : CascadeMux
    port map (
            O => \N__34560\,
            I => \N__34557\
        );

    \I__6923\ : InMux
    port map (
            O => \N__34557\,
            I => \N__34554\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__34554\,
            I => \N__34551\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__34551\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__34548\,
            I => \N__34545\
        );

    \I__6919\ : InMux
    port map (
            O => \N__34545\,
            I => \N__34542\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__34542\,
            I => \N__34539\
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__34539\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__6916\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34533\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__34533\,
            I => \N__34530\
        );

    \I__6914\ : Odrv4
    port map (
            O => \N__34530\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__34527\,
            I => \N__34524\
        );

    \I__6912\ : InMux
    port map (
            O => \N__34524\,
            I => \N__34521\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__34521\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__6910\ : InMux
    port map (
            O => \N__34518\,
            I => \N__34515\
        );

    \I__6909\ : LocalMux
    port map (
            O => \N__34515\,
            I => \N__34512\
        );

    \I__6908\ : Span4Mux_h
    port map (
            O => \N__34512\,
            I => \N__34509\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__34509\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__6906\ : CascadeMux
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__6905\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34500\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__34500\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__6903\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34494\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__34494\,
            I => \N__34491\
        );

    \I__6901\ : Odrv12
    port map (
            O => \N__34491\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__6900\ : CascadeMux
    port map (
            O => \N__34488\,
            I => \N__34485\
        );

    \I__6899\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34482\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__34482\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__34479\,
            I => \N__34476\
        );

    \I__6896\ : InMux
    port map (
            O => \N__34476\,
            I => \N__34473\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34470\
        );

    \I__6894\ : Odrv4
    port map (
            O => \N__34470\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__6893\ : InMux
    port map (
            O => \N__34467\,
            I => \N__34464\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__34464\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__6891\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34458\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__34458\,
            I => \N__34455\
        );

    \I__6889\ : Odrv4
    port map (
            O => \N__34455\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__34452\,
            I => \N__34449\
        );

    \I__6887\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34446\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__6885\ : Odrv4
    port map (
            O => \N__34443\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__6884\ : InMux
    port map (
            O => \N__34440\,
            I => \N__34437\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34437\,
            I => \N__34434\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__34434\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__34431\,
            I => \N__34428\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34425\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34425\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__6878\ : CascadeMux
    port map (
            O => \N__34422\,
            I => \N__34419\
        );

    \I__6877\ : InMux
    port map (
            O => \N__34419\,
            I => \N__34416\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34416\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__6875\ : InMux
    port map (
            O => \N__34413\,
            I => \N__34410\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__34410\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__6873\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34404\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__34404\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34398\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__34398\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__6869\ : CascadeMux
    port map (
            O => \N__34395\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\
        );

    \I__6868\ : CascadeMux
    port map (
            O => \N__34392\,
            I => \N__34389\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34389\,
            I => \N__34386\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__34386\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34380\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__34380\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34371\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34371\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__34368\,
            I => \N__34365\
        );

    \I__6859\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34362\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__34362\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__6857\ : CascadeMux
    port map (
            O => \N__34359\,
            I => \N__34356\
        );

    \I__6856\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__34353\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__6854\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34322\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34322\
        );

    \I__6852\ : InMux
    port map (
            O => \N__34348\,
            I => \N__34322\
        );

    \I__6851\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34322\
        );

    \I__6850\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34313\
        );

    \I__6849\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34313\
        );

    \I__6848\ : InMux
    port map (
            O => \N__34344\,
            I => \N__34313\
        );

    \I__6847\ : InMux
    port map (
            O => \N__34343\,
            I => \N__34313\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34342\,
            I => \N__34294\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34341\,
            I => \N__34294\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34340\,
            I => \N__34294\
        );

    \I__6843\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34294\
        );

    \I__6842\ : InMux
    port map (
            O => \N__34338\,
            I => \N__34285\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34337\,
            I => \N__34285\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34336\,
            I => \N__34285\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34285\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34276\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34276\
        );

    \I__6836\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34276\
        );

    \I__6835\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34276\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34271\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__34313\,
            I => \N__34271\
        );

    \I__6832\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34266\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34311\,
            I => \N__34266\
        );

    \I__6830\ : InMux
    port map (
            O => \N__34310\,
            I => \N__34257\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34257\
        );

    \I__6828\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34257\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34307\,
            I => \N__34257\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34248\
        );

    \I__6825\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34248\
        );

    \I__6824\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34248\
        );

    \I__6823\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34248\
        );

    \I__6822\ : LocalMux
    port map (
            O => \N__34294\,
            I => \N__34245\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__34285\,
            I => \N__34238\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34238\
        );

    \I__6819\ : Span4Mux_h
    port map (
            O => \N__34271\,
            I => \N__34238\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__34266\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__34257\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__34248\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6815\ : Odrv12
    port map (
            O => \N__34245\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__34238\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__34227\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__34221\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__6810\ : CascadeMux
    port map (
            O => \N__34218\,
            I => \N__34214\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__34217\,
            I => \N__34211\
        );

    \I__6808\ : InMux
    port map (
            O => \N__34214\,
            I => \N__34205\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34211\,
            I => \N__34205\
        );

    \I__6806\ : InMux
    port map (
            O => \N__34210\,
            I => \N__34202\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__34205\,
            I => \N__34199\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6803\ : Odrv4
    port map (
            O => \N__34199\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34194\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34184\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34184\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34181\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__34184\,
            I => \N__34178\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__34181\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6796\ : Odrv4
    port map (
            O => \N__34178\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34173\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__6794\ : CascadeMux
    port map (
            O => \N__34170\,
            I => \N__34166\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34163\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34159\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34163\,
            I => \N__34156\
        );

    \I__6790\ : InMux
    port map (
            O => \N__34162\,
            I => \N__34153\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__34159\,
            I => \N__34148\
        );

    \I__6788\ : Span4Mux_h
    port map (
            O => \N__34156\,
            I => \N__34148\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34153\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6786\ : Odrv4
    port map (
            O => \N__34148\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__6785\ : InMux
    port map (
            O => \N__34143\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34140\,
            I => \N__34136\
        );

    \I__6783\ : CascadeMux
    port map (
            O => \N__34139\,
            I => \N__34132\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34136\,
            I => \N__34129\
        );

    \I__6781\ : InMux
    port map (
            O => \N__34135\,
            I => \N__34126\
        );

    \I__6780\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34123\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__34129\,
            I => \N__34120\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__34126\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__34123\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6776\ : Odrv4
    port map (
            O => \N__34120\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__6775\ : InMux
    port map (
            O => \N__34113\,
            I => \bfn_14_8_0_\
        );

    \I__6774\ : CascadeMux
    port map (
            O => \N__34110\,
            I => \N__34107\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34104\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__34104\,
            I => \N__34100\
        );

    \I__6771\ : InMux
    port map (
            O => \N__34103\,
            I => \N__34096\
        );

    \I__6770\ : Span4Mux_h
    port map (
            O => \N__34100\,
            I => \N__34093\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34099\,
            I => \N__34090\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__34096\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__34093\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__34090\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34083\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__6764\ : CascadeMux
    port map (
            O => \N__34080\,
            I => \N__34076\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__34079\,
            I => \N__34073\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34076\,
            I => \N__34067\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34067\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34072\,
            I => \N__34064\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__34067\,
            I => \N__34061\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__34064\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6757\ : Odrv4
    port map (
            O => \N__34061\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34056\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34053\,
            I => \N__34046\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34052\,
            I => \N__34046\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34043\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__34040\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__34043\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__34040\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34035\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__6748\ : InMux
    port map (
            O => \N__34032\,
            I => \N__34028\
        );

    \I__6747\ : InMux
    port map (
            O => \N__34031\,
            I => \N__34025\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__34028\,
            I => \N__34022\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__34025\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6744\ : Odrv4
    port map (
            O => \N__34022\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34017\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34014\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__6741\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \N__34008\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34004\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34007\,
            I => \N__34001\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34004\,
            I => \N__33998\
        );

    \I__6737\ : LocalMux
    port map (
            O => \N__34001\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__33998\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__6735\ : CEMux
    port map (
            O => \N__33993\,
            I => \N__33988\
        );

    \I__6734\ : CEMux
    port map (
            O => \N__33992\,
            I => \N__33985\
        );

    \I__6733\ : CEMux
    port map (
            O => \N__33991\,
            I => \N__33981\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__33988\,
            I => \N__33978\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__33985\,
            I => \N__33975\
        );

    \I__6730\ : CEMux
    port map (
            O => \N__33984\,
            I => \N__33972\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__33981\,
            I => \N__33969\
        );

    \I__6728\ : Span4Mux_v
    port map (
            O => \N__33978\,
            I => \N__33962\
        );

    \I__6727\ : Span4Mux_v
    port map (
            O => \N__33975\,
            I => \N__33962\
        );

    \I__6726\ : LocalMux
    port map (
            O => \N__33972\,
            I => \N__33962\
        );

    \I__6725\ : Span4Mux_v
    port map (
            O => \N__33969\,
            I => \N__33959\
        );

    \I__6724\ : Span4Mux_v
    port map (
            O => \N__33962\,
            I => \N__33956\
        );

    \I__6723\ : Span4Mux_v
    port map (
            O => \N__33959\,
            I => \N__33953\
        );

    \I__6722\ : Span4Mux_v
    port map (
            O => \N__33956\,
            I => \N__33950\
        );

    \I__6721\ : Span4Mux_v
    port map (
            O => \N__33953\,
            I => \N__33947\
        );

    \I__6720\ : Span4Mux_v
    port map (
            O => \N__33950\,
            I => \N__33944\
        );

    \I__6719\ : Odrv4
    port map (
            O => \N__33947\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__33944\,
            I => \delay_measurement_inst.delay_tr_timer.N_201_i\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__33939\,
            I => \N__33935\
        );

    \I__6716\ : CascadeMux
    port map (
            O => \N__33938\,
            I => \N__33932\
        );

    \I__6715\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33926\
        );

    \I__6714\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33926\
        );

    \I__6713\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33923\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__33926\,
            I => \N__33920\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__33923\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6710\ : Odrv4
    port map (
            O => \N__33920\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__6709\ : InMux
    port map (
            O => \N__33915\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__33912\,
            I => \N__33908\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__33911\,
            I => \N__33905\
        );

    \I__6706\ : InMux
    port map (
            O => \N__33908\,
            I => \N__33900\
        );

    \I__6705\ : InMux
    port map (
            O => \N__33905\,
            I => \N__33900\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__33900\,
            I => \N__33896\
        );

    \I__6703\ : InMux
    port map (
            O => \N__33899\,
            I => \N__33893\
        );

    \I__6702\ : Span4Mux_h
    port map (
            O => \N__33896\,
            I => \N__33890\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__33893\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6700\ : Odrv4
    port map (
            O => \N__33890\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__6699\ : InMux
    port map (
            O => \N__33885\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__33882\,
            I => \N__33878\
        );

    \I__6697\ : InMux
    port map (
            O => \N__33881\,
            I => \N__33875\
        );

    \I__6696\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33871\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__33875\,
            I => \N__33868\
        );

    \I__6694\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33865\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33860\
        );

    \I__6692\ : Span4Mux_h
    port map (
            O => \N__33868\,
            I => \N__33860\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__33865\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__33860\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__6689\ : InMux
    port map (
            O => \N__33855\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__33852\,
            I => \N__33849\
        );

    \I__6687\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__33846\,
            I => \N__33841\
        );

    \I__6685\ : InMux
    port map (
            O => \N__33845\,
            I => \N__33838\
        );

    \I__6684\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33835\
        );

    \I__6683\ : Odrv4
    port map (
            O => \N__33841\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__33838\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__33835\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__6680\ : InMux
    port map (
            O => \N__33828\,
            I => \bfn_14_7_0_\
        );

    \I__6679\ : CascadeMux
    port map (
            O => \N__33825\,
            I => \N__33822\
        );

    \I__6678\ : InMux
    port map (
            O => \N__33822\,
            I => \N__33819\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__33819\,
            I => \N__33815\
        );

    \I__6676\ : InMux
    port map (
            O => \N__33818\,
            I => \N__33811\
        );

    \I__6675\ : Span4Mux_h
    port map (
            O => \N__33815\,
            I => \N__33808\
        );

    \I__6674\ : InMux
    port map (
            O => \N__33814\,
            I => \N__33805\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__33811\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__33808\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6671\ : LocalMux
    port map (
            O => \N__33805\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__6670\ : InMux
    port map (
            O => \N__33798\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__6669\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33788\
        );

    \I__6668\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33788\
        );

    \I__6667\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33785\
        );

    \I__6666\ : LocalMux
    port map (
            O => \N__33788\,
            I => \N__33782\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33777\
        );

    \I__6664\ : Span4Mux_v
    port map (
            O => \N__33782\,
            I => \N__33777\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__33777\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__6662\ : InMux
    port map (
            O => \N__33774\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__6661\ : InMux
    port map (
            O => \N__33771\,
            I => \N__33764\
        );

    \I__6660\ : InMux
    port map (
            O => \N__33770\,
            I => \N__33764\
        );

    \I__6659\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33761\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__33764\,
            I => \N__33758\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__33761\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__33758\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__6655\ : InMux
    port map (
            O => \N__33753\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__33750\,
            I => \N__33746\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__33749\,
            I => \N__33743\
        );

    \I__6652\ : InMux
    port map (
            O => \N__33746\,
            I => \N__33738\
        );

    \I__6651\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33738\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33734\
        );

    \I__6649\ : InMux
    port map (
            O => \N__33737\,
            I => \N__33731\
        );

    \I__6648\ : Span4Mux_h
    port map (
            O => \N__33734\,
            I => \N__33728\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__33731\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6646\ : Odrv4
    port map (
            O => \N__33728\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__6645\ : InMux
    port map (
            O => \N__33723\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__33720\,
            I => \N__33716\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__33719\,
            I => \N__33713\
        );

    \I__6642\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33707\
        );

    \I__6641\ : InMux
    port map (
            O => \N__33713\,
            I => \N__33707\
        );

    \I__6640\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33704\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__33707\,
            I => \N__33701\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__33704\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6637\ : Odrv4
    port map (
            O => \N__33701\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__6636\ : InMux
    port map (
            O => \N__33696\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__6635\ : CascadeMux
    port map (
            O => \N__33693\,
            I => \N__33689\
        );

    \I__6634\ : CascadeMux
    port map (
            O => \N__33692\,
            I => \N__33686\
        );

    \I__6633\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33681\
        );

    \I__6632\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33681\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__33681\,
            I => \N__33677\
        );

    \I__6630\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33674\
        );

    \I__6629\ : Span4Mux_h
    port map (
            O => \N__33677\,
            I => \N__33671\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__33674\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__33671\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__6626\ : InMux
    port map (
            O => \N__33666\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__6625\ : CascadeMux
    port map (
            O => \N__33663\,
            I => \N__33660\
        );

    \I__6624\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33656\
        );

    \I__6623\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33653\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__33656\,
            I => \N__33647\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33647\
        );

    \I__6620\ : InMux
    port map (
            O => \N__33652\,
            I => \N__33644\
        );

    \I__6619\ : Span4Mux_h
    port map (
            O => \N__33647\,
            I => \N__33641\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__33644\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__33641\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__6616\ : InMux
    port map (
            O => \N__33636\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__6615\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33630\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__6613\ : Span4Mux_h
    port map (
            O => \N__33627\,
            I => \N__33622\
        );

    \I__6612\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33619\
        );

    \I__6611\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33616\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__33622\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__33619\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__33616\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__6607\ : InMux
    port map (
            O => \N__33609\,
            I => \bfn_14_6_0_\
        );

    \I__6606\ : CascadeMux
    port map (
            O => \N__33606\,
            I => \N__33603\
        );

    \I__6605\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33600\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__33600\,
            I => \N__33596\
        );

    \I__6603\ : InMux
    port map (
            O => \N__33599\,
            I => \N__33592\
        );

    \I__6602\ : Span4Mux_h
    port map (
            O => \N__33596\,
            I => \N__33589\
        );

    \I__6601\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33586\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__33592\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6599\ : Odrv4
    port map (
            O => \N__33589\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__33586\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__6597\ : InMux
    port map (
            O => \N__33579\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__33576\,
            I => \N__33572\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__33575\,
            I => \N__33569\
        );

    \I__6594\ : InMux
    port map (
            O => \N__33572\,
            I => \N__33563\
        );

    \I__6593\ : InMux
    port map (
            O => \N__33569\,
            I => \N__33563\
        );

    \I__6592\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33560\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__33563\,
            I => \N__33557\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__33560\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6589\ : Odrv4
    port map (
            O => \N__33557\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__6588\ : InMux
    port map (
            O => \N__33552\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__6587\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33542\
        );

    \I__6586\ : InMux
    port map (
            O => \N__33548\,
            I => \N__33542\
        );

    \I__6585\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33539\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__33542\,
            I => \N__33536\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__33539\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__33536\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__6581\ : InMux
    port map (
            O => \N__33531\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__6580\ : InMux
    port map (
            O => \N__33528\,
            I => \N__33521\
        );

    \I__6579\ : InMux
    port map (
            O => \N__33527\,
            I => \N__33521\
        );

    \I__6578\ : InMux
    port map (
            O => \N__33526\,
            I => \N__33518\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__33521\,
            I => \N__33515\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__33518\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6575\ : Odrv4
    port map (
            O => \N__33515\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__6574\ : InMux
    port map (
            O => \N__33510\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__6573\ : CascadeMux
    port map (
            O => \N__33507\,
            I => \N__33504\
        );

    \I__6572\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__33501\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__6570\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__33495\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__6568\ : InMux
    port map (
            O => \N__33492\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__6567\ : IoInMux
    port map (
            O => \N__33489\,
            I => \N__33486\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__6565\ : Span4Mux_s2_v
    port map (
            O => \N__33483\,
            I => \N__33480\
        );

    \I__6564\ : Sp12to4
    port map (
            O => \N__33480\,
            I => \N__33477\
        );

    \I__6563\ : Span12Mux_h
    port map (
            O => \N__33477\,
            I => \N__33474\
        );

    \I__6562\ : Span12Mux_v
    port map (
            O => \N__33474\,
            I => \N__33471\
        );

    \I__6561\ : Odrv12
    port map (
            O => \N__33471\,
            I => pwm_output_c
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__33468\,
            I => \N__33465\
        );

    \I__6559\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33462\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__33462\,
            I => \N__33458\
        );

    \I__6557\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33454\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__33458\,
            I => \N__33450\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33457\,
            I => \N__33447\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__33454\,
            I => \N__33444\
        );

    \I__6553\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33441\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__33450\,
            I => \N__33438\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__33447\,
            I => \N__33433\
        );

    \I__6550\ : Span12Mux_v
    port map (
            O => \N__33444\,
            I => \N__33433\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__33441\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6548\ : Odrv4
    port map (
            O => \N__33438\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__33433\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6546\ : IoInMux
    port map (
            O => \N__33426\,
            I => \N__33423\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__33423\,
            I => \N__33420\
        );

    \I__6544\ : Odrv4
    port map (
            O => \N__33420\,
            I => s2_phy_c
        );

    \I__6543\ : InMux
    port map (
            O => \N__33417\,
            I => \bfn_14_5_0_\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__33414\,
            I => \N__33411\
        );

    \I__6541\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33408\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33403\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33400\
        );

    \I__6538\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33397\
        );

    \I__6537\ : Span4Mux_h
    port map (
            O => \N__33403\,
            I => \N__33394\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__33400\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__33397\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6534\ : Odrv4
    port map (
            O => \N__33394\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33387\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__6531\ : InMux
    port map (
            O => \N__33381\,
            I => \N__33376\
        );

    \I__6530\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33373\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33370\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__33376\,
            I => \N__33365\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33365\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33360\
        );

    \I__6525\ : Span4Mux_v
    port map (
            O => \N__33365\,
            I => \N__33360\
        );

    \I__6524\ : Odrv4
    port map (
            O => \N__33360\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33357\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__6522\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33347\
        );

    \I__6521\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33347\
        );

    \I__6520\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33344\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__33347\,
            I => \N__33341\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33344\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__33341\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__6516\ : InMux
    port map (
            O => \N__33336\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33333\,
            I => \N__33326\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33332\,
            I => \N__33326\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33323\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__33326\,
            I => \N__33320\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__33323\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__33320\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33315\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__6508\ : CascadeMux
    port map (
            O => \N__33312\,
            I => \N__33309\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33309\,
            I => \N__33306\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__33306\,
            I => \pwm_generator_inst.un14_counter_1\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33300\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__6502\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33291\
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__6500\ : Odrv12
    port map (
            O => \N__33288\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__6499\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33282\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__33282\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__6497\ : CascadeMux
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33276\,
            I => \N__33273\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__33273\,
            I => \N__33270\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__33270\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__6493\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33264\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33264\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33258\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33258\,
            I => \N__33255\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33252\
        );

    \I__6488\ : Odrv12
    port map (
            O => \N__33252\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__6487\ : InMux
    port map (
            O => \N__33249\,
            I => \N__33246\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__33246\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__33243\,
            I => \N__33240\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33237\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__33237\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33231\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__33231\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__33228\,
            I => \N__33225\
        );

    \I__6479\ : InMux
    port map (
            O => \N__33225\,
            I => \N__33222\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33222\,
            I => \pwm_generator_inst.un14_counter_6\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33219\,
            I => \N__33216\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__33216\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__6475\ : CascadeMux
    port map (
            O => \N__33213\,
            I => \N__33210\
        );

    \I__6474\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__33207\,
            I => \pwm_generator_inst.un14_counter_7\
        );

    \I__6472\ : InMux
    port map (
            O => \N__33204\,
            I => \N__33201\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33201\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__33198\,
            I => \N__33195\
        );

    \I__6469\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__33192\,
            I => \N__33189\
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__33189\,
            I => \pwm_generator_inst.un14_counter_8\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33186\,
            I => \N__33183\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__33183\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33180\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33177\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33174\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33171\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33168\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33165\,
            I => \bfn_13_23_0_\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33162\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33156\
        );

    \I__6456\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33152\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33148\
        );

    \I__6454\ : Span12Mux_v
    port map (
            O => \N__33152\,
            I => \N__33145\
        );

    \I__6453\ : InMux
    port map (
            O => \N__33151\,
            I => \N__33142\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33148\,
            I => \N__33139\
        );

    \I__6451\ : Odrv12
    port map (
            O => \N__33145\,
            I => \il_min_comp1_D2\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__33142\,
            I => \il_min_comp1_D2\
        );

    \I__6449\ : Odrv12
    port map (
            O => \N__33139\,
            I => \il_min_comp1_D2\
        );

    \I__6448\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33128\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33125\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__33128\,
            I => \N__33122\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33119\
        );

    \I__6444\ : Span4Mux_v
    port map (
            O => \N__33122\,
            I => \N__33116\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__33119\,
            I => \N__33113\
        );

    \I__6442\ : Span4Mux_v
    port map (
            O => \N__33116\,
            I => \N__33110\
        );

    \I__6441\ : Span12Mux_s7_v
    port map (
            O => \N__33113\,
            I => \N__33107\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__33110\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__6439\ : Odrv12
    port map (
            O => \N__33107\,
            I => \phase_controller_inst1.state_RNIE87FZ0Z_2\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__33099\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__6436\ : InMux
    port map (
            O => \N__33096\,
            I => \N__33093\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__33093\,
            I => \N__33090\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__33090\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33083\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33080\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33083\,
            I => \N__33073\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33080\,
            I => \N__33073\
        );

    \I__6429\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33070\
        );

    \I__6428\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33067\
        );

    \I__6427\ : Odrv12
    port map (
            O => \N__33073\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__33070\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__33067\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__6424\ : CascadeMux
    port map (
            O => \N__33060\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__6423\ : CascadeMux
    port map (
            O => \N__33057\,
            I => \N__33054\
        );

    \I__6422\ : InMux
    port map (
            O => \N__33054\,
            I => \N__33051\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__33051\,
            I => \N__33048\
        );

    \I__6420\ : Span4Mux_h
    port map (
            O => \N__33048\,
            I => \N__33045\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__33045\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33042\,
            I => \N__33032\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33041\,
            I => \N__33032\
        );

    \I__6416\ : InMux
    port map (
            O => \N__33040\,
            I => \N__33032\
        );

    \I__6415\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33029\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__33032\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__33029\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6412\ : CascadeMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__6411\ : InMux
    port map (
            O => \N__33021\,
            I => \N__33013\
        );

    \I__6410\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33013\
        );

    \I__6409\ : InMux
    port map (
            O => \N__33019\,
            I => \N__33010\
        );

    \I__6408\ : InMux
    port map (
            O => \N__33018\,
            I => \N__33007\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__33013\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33010\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__33007\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6404\ : IoInMux
    port map (
            O => \N__33000\,
            I => \N__32997\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__32997\,
            I => \N__32994\
        );

    \I__6402\ : Odrv12
    port map (
            O => \N__32994\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__6401\ : InMux
    port map (
            O => \N__32991\,
            I => \bfn_13_22_0_\
        );

    \I__6400\ : InMux
    port map (
            O => \N__32988\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__6399\ : InMux
    port map (
            O => \N__32985\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__6398\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32979\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__32979\,
            I => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\
        );

    \I__6396\ : CascadeMux
    port map (
            O => \N__32976\,
            I => \N__32973\
        );

    \I__6395\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32970\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__32970\,
            I => \N__32967\
        );

    \I__6393\ : Odrv4
    port map (
            O => \N__32967\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__6392\ : InMux
    port map (
            O => \N__32964\,
            I => \N__32961\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__32961\,
            I => \N__32958\
        );

    \I__6390\ : Span4Mux_h
    port map (
            O => \N__32958\,
            I => \N__32955\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__32955\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__32952\,
            I => \N__32949\
        );

    \I__6387\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32946\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__32946\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__6385\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32940\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__6383\ : Odrv4
    port map (
            O => \N__32937\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__6382\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__32931\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__32928\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\
        );

    \I__6379\ : InMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32918\
        );

    \I__6377\ : InMux
    port map (
            O => \N__32921\,
            I => \N__32915\
        );

    \I__6376\ : Odrv12
    port map (
            O => \N__32918\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__32915\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__6374\ : InMux
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__32907\,
            I => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\
        );

    \I__6372\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32901\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__32901\,
            I => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\
        );

    \I__6370\ : InMux
    port map (
            O => \N__32898\,
            I => \N__32895\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__32895\,
            I => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\
        );

    \I__6368\ : CascadeMux
    port map (
            O => \N__32892\,
            I => \N__32888\
        );

    \I__6367\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32885\
        );

    \I__6366\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32882\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__32885\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__32882\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__6363\ : InMux
    port map (
            O => \N__32877\,
            I => \N__32874\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__32874\,
            I => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\
        );

    \I__6361\ : CascadeMux
    port map (
            O => \N__32871\,
            I => \N__32868\
        );

    \I__6360\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32865\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__32865\,
            I => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\
        );

    \I__6358\ : InMux
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__32859\,
            I => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__32856\,
            I => \N__32853\
        );

    \I__6355\ : InMux
    port map (
            O => \N__32853\,
            I => \N__32850\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__32850\,
            I => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\
        );

    \I__6353\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32844\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__32844\,
            I => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__32841\,
            I => \N__32838\
        );

    \I__6350\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32835\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__32835\,
            I => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\
        );

    \I__6348\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32829\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__32829\,
            I => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\
        );

    \I__6346\ : CascadeMux
    port map (
            O => \N__32826\,
            I => \N__32823\
        );

    \I__6345\ : InMux
    port map (
            O => \N__32823\,
            I => \N__32820\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__32820\,
            I => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\
        );

    \I__6343\ : CascadeMux
    port map (
            O => \N__32817\,
            I => \N__32814\
        );

    \I__6342\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32811\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__32811\,
            I => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__32808\,
            I => \N__32804\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__32807\,
            I => \N__32801\
        );

    \I__6338\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32798\
        );

    \I__6337\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32793\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__32798\,
            I => \N__32790\
        );

    \I__6335\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32787\
        );

    \I__6334\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32784\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__32793\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__32790\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__32787\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__32784\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__32775\,
            I => \N__32772\
        );

    \I__6328\ : InMux
    port map (
            O => \N__32772\,
            I => \N__32769\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__32769\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__6326\ : InMux
    port map (
            O => \N__32766\,
            I => \N__32763\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__32763\,
            I => \N__32760\
        );

    \I__6324\ : Span4Mux_v
    port map (
            O => \N__32760\,
            I => \N__32757\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__32757\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__32754\,
            I => \N__32750\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__32753\,
            I => \N__32746\
        );

    \I__6320\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32741\
        );

    \I__6319\ : InMux
    port map (
            O => \N__32749\,
            I => \N__32741\
        );

    \I__6318\ : InMux
    port map (
            O => \N__32746\,
            I => \N__32738\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__32741\,
            I => \N__32735\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__32738\,
            I => \N__32732\
        );

    \I__6315\ : Span4Mux_v
    port map (
            O => \N__32735\,
            I => \N__32726\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__32732\,
            I => \N__32726\
        );

    \I__6313\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32723\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__32726\,
            I => \N__32720\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__32723\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__32720\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6309\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32710\
        );

    \I__6308\ : InMux
    port map (
            O => \N__32714\,
            I => \N__32705\
        );

    \I__6307\ : InMux
    port map (
            O => \N__32713\,
            I => \N__32705\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__32710\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__32705\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6304\ : InMux
    port map (
            O => \N__32700\,
            I => \N__32696\
        );

    \I__6303\ : InMux
    port map (
            O => \N__32699\,
            I => \N__32693\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__32696\,
            I => \N__32690\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__32693\,
            I => \N__32684\
        );

    \I__6300\ : Span4Mux_v
    port map (
            O => \N__32690\,
            I => \N__32684\
        );

    \I__6299\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32681\
        );

    \I__6298\ : Sp12to4
    port map (
            O => \N__32684\,
            I => \N__32678\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__32681\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6296\ : Odrv12
    port map (
            O => \N__32678\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6295\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32669\
        );

    \I__6294\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32666\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__32669\,
            I => \N__32661\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__32666\,
            I => \N__32661\
        );

    \I__6291\ : Span4Mux_s3_v
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__6290\ : Span4Mux_h
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__6289\ : Sp12to4
    port map (
            O => \N__32655\,
            I => \N__32650\
        );

    \I__6288\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32645\
        );

    \I__6287\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32645\
        );

    \I__6286\ : Span12Mux_v
    port map (
            O => \N__32650\,
            I => \N__32642\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__32645\,
            I => \N__32639\
        );

    \I__6284\ : Span12Mux_v
    port map (
            O => \N__32642\,
            I => \N__32636\
        );

    \I__6283\ : Span12Mux_h
    port map (
            O => \N__32639\,
            I => \N__32633\
        );

    \I__6282\ : Span12Mux_h
    port map (
            O => \N__32636\,
            I => \N__32628\
        );

    \I__6281\ : Span12Mux_v
    port map (
            O => \N__32633\,
            I => \N__32628\
        );

    \I__6280\ : Odrv12
    port map (
            O => \N__32628\,
            I => start_stop_c
        );

    \I__6279\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32622\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__32622\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__6277\ : CascadeMux
    port map (
            O => \N__32619\,
            I => \N__32616\
        );

    \I__6276\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32610\
        );

    \I__6275\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32610\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__32610\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__6273\ : CascadeMux
    port map (
            O => \N__32607\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\
        );

    \I__6272\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32598\
        );

    \I__6271\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32598\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__32598\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__32595\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\
        );

    \I__6268\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32583\
        );

    \I__6267\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32583\
        );

    \I__6266\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32583\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__32583\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__6264\ : InMux
    port map (
            O => \N__32580\,
            I => \N__32571\
        );

    \I__6263\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32571\
        );

    \I__6262\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32571\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__32571\,
            I => \N__32568\
        );

    \I__6260\ : Span4Mux_v
    port map (
            O => \N__32568\,
            I => \N__32565\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__32565\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__6258\ : InMux
    port map (
            O => \N__32562\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__6257\ : InMux
    port map (
            O => \N__32559\,
            I => \bfn_13_10_0_\
        );

    \I__6256\ : InMux
    port map (
            O => \N__32556\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__6255\ : InMux
    port map (
            O => \N__32553\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__6254\ : InMux
    port map (
            O => \N__32550\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__6253\ : InMux
    port map (
            O => \N__32547\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__6252\ : CascadeMux
    port map (
            O => \N__32544\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\
        );

    \I__6251\ : InMux
    port map (
            O => \N__32541\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__6250\ : InMux
    port map (
            O => \N__32538\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__6249\ : InMux
    port map (
            O => \N__32535\,
            I => \bfn_13_9_0_\
        );

    \I__6248\ : InMux
    port map (
            O => \N__32532\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__6247\ : InMux
    port map (
            O => \N__32529\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__6246\ : InMux
    port map (
            O => \N__32526\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__6245\ : InMux
    port map (
            O => \N__32523\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__6244\ : InMux
    port map (
            O => \N__32520\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__6243\ : InMux
    port map (
            O => \N__32517\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__6242\ : InMux
    port map (
            O => \N__32514\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__6241\ : InMux
    port map (
            O => \N__32511\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__6240\ : InMux
    port map (
            O => \N__32508\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__6239\ : InMux
    port map (
            O => \N__32505\,
            I => \bfn_13_8_0_\
        );

    \I__6238\ : InMux
    port map (
            O => \N__32502\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__6237\ : InMux
    port map (
            O => \N__32499\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__6236\ : InMux
    port map (
            O => \N__32496\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__6235\ : InMux
    port map (
            O => \N__32493\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__6234\ : InMux
    port map (
            O => \N__32490\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__6233\ : IoInMux
    port map (
            O => \N__32487\,
            I => \N__32484\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__32484\,
            I => \N__32481\
        );

    \I__6231\ : Span4Mux_s0_v
    port map (
            O => \N__32481\,
            I => \N__32471\
        );

    \I__6230\ : InMux
    port map (
            O => \N__32480\,
            I => \N__32440\
        );

    \I__6229\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32440\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32478\,
            I => \N__32440\
        );

    \I__6227\ : InMux
    port map (
            O => \N__32477\,
            I => \N__32431\
        );

    \I__6226\ : InMux
    port map (
            O => \N__32476\,
            I => \N__32431\
        );

    \I__6225\ : InMux
    port map (
            O => \N__32475\,
            I => \N__32431\
        );

    \I__6224\ : InMux
    port map (
            O => \N__32474\,
            I => \N__32431\
        );

    \I__6223\ : Sp12to4
    port map (
            O => \N__32471\,
            I => \N__32428\
        );

    \I__6222\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32425\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32416\
        );

    \I__6220\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32416\
        );

    \I__6219\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32416\
        );

    \I__6218\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32416\
        );

    \I__6217\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32407\
        );

    \I__6216\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32407\
        );

    \I__6215\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32407\
        );

    \I__6214\ : InMux
    port map (
            O => \N__32462\,
            I => \N__32407\
        );

    \I__6213\ : InMux
    port map (
            O => \N__32461\,
            I => \N__32400\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32460\,
            I => \N__32400\
        );

    \I__6211\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32400\
        );

    \I__6210\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32391\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32391\
        );

    \I__6208\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32391\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32391\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32382\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32453\,
            I => \N__32382\
        );

    \I__6204\ : InMux
    port map (
            O => \N__32452\,
            I => \N__32382\
        );

    \I__6203\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32382\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32450\,
            I => \N__32373\
        );

    \I__6201\ : InMux
    port map (
            O => \N__32449\,
            I => \N__32373\
        );

    \I__6200\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32373\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32447\,
            I => \N__32373\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__32440\,
            I => \N__32368\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__32431\,
            I => \N__32368\
        );

    \I__6196\ : Span12Mux_s5_h
    port map (
            O => \N__32428\,
            I => \N__32365\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__32425\,
            I => \N__32362\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32416\,
            I => \N__32357\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32357\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__32400\,
            I => \N__32348\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__32391\,
            I => \N__32348\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__32382\,
            I => \N__32348\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32373\,
            I => \N__32348\
        );

    \I__6188\ : Span4Mux_h
    port map (
            O => \N__32368\,
            I => \N__32345\
        );

    \I__6187\ : Span12Mux_v
    port map (
            O => \N__32365\,
            I => \N__32342\
        );

    \I__6186\ : Span12Mux_h
    port map (
            O => \N__32362\,
            I => \N__32339\
        );

    \I__6185\ : Span4Mux_v
    port map (
            O => \N__32357\,
            I => \N__32334\
        );

    \I__6184\ : Span4Mux_v
    port map (
            O => \N__32348\,
            I => \N__32334\
        );

    \I__6183\ : Span4Mux_v
    port map (
            O => \N__32345\,
            I => \N__32331\
        );

    \I__6182\ : Span12Mux_v
    port map (
            O => \N__32342\,
            I => \N__32328\
        );

    \I__6181\ : Odrv12
    port map (
            O => \N__32339\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6180\ : Odrv4
    port map (
            O => \N__32334\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__32331\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6178\ : Odrv12
    port map (
            O => \N__32328\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__6177\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32316\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__32316\,
            I => \N__32312\
        );

    \I__6175\ : CascadeMux
    port map (
            O => \N__32315\,
            I => \N__32309\
        );

    \I__6174\ : Span4Mux_h
    port map (
            O => \N__32312\,
            I => \N__32306\
        );

    \I__6173\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32303\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__32306\,
            I => \N__32300\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32303\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__32300\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__6169\ : CascadeMux
    port map (
            O => \N__32295\,
            I => \N__32291\
        );

    \I__6168\ : InMux
    port map (
            O => \N__32294\,
            I => \N__32280\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32291\,
            I => \N__32280\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32290\,
            I => \N__32280\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32289\,
            I => \N__32280\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__32280\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__6163\ : InMux
    port map (
            O => \N__32277\,
            I => \N__32265\
        );

    \I__6162\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32265\
        );

    \I__6161\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32265\
        );

    \I__6160\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32265\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32262\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__32262\,
            I => \N__32259\
        );

    \I__6157\ : Odrv4
    port map (
            O => \N__32259\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32256\,
            I => \N__32253\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32253\,
            I => \N__32250\
        );

    \I__6154\ : Span4Mux_h
    port map (
            O => \N__32250\,
            I => \N__32246\
        );

    \I__6153\ : InMux
    port map (
            O => \N__32249\,
            I => \N__32243\
        );

    \I__6152\ : Span4Mux_v
    port map (
            O => \N__32246\,
            I => \N__32240\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32243\,
            I => \N__32237\
        );

    \I__6150\ : Odrv4
    port map (
            O => \N__32240\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__6149\ : Odrv12
    port map (
            O => \N__32237\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__6148\ : CascadeMux
    port map (
            O => \N__32232\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32229\,
            I => \N__32225\
        );

    \I__6146\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32222\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__32225\,
            I => \N__32217\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32222\,
            I => \N__32217\
        );

    \I__6143\ : Span4Mux_v
    port map (
            O => \N__32217\,
            I => \N__32211\
        );

    \I__6142\ : InMux
    port map (
            O => \N__32216\,
            I => \N__32204\
        );

    \I__6141\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32204\
        );

    \I__6140\ : InMux
    port map (
            O => \N__32214\,
            I => \N__32204\
        );

    \I__6139\ : Odrv4
    port map (
            O => \N__32211\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__32204\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__6137\ : InMux
    port map (
            O => \N__32199\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32196\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32193\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__6134\ : InMux
    port map (
            O => \N__32190\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__6133\ : InMux
    port map (
            O => \N__32187\,
            I => \N__32184\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32184\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__6131\ : CascadeMux
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__6130\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32175\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__32175\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\
        );

    \I__6128\ : IoInMux
    port map (
            O => \N__32172\,
            I => \N__32169\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32169\,
            I => \N__32166\
        );

    \I__6126\ : Span4Mux_s0_v
    port map (
            O => \N__32166\,
            I => \N__32163\
        );

    \I__6125\ : Odrv4
    port map (
            O => \N__32163\,
            I => \pll_inst.red_c_i\
        );

    \I__6124\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32154\
        );

    \I__6123\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32147\
        );

    \I__6122\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32147\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32147\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__32154\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__32147\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6118\ : CascadeMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32134\
        );

    \I__6116\ : InMux
    port map (
            O => \N__32138\,
            I => \N__32129\
        );

    \I__6115\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32129\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__32134\,
            I => \N__32126\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32123\
        );

    \I__6112\ : Span4Mux_h
    port map (
            O => \N__32126\,
            I => \N__32120\
        );

    \I__6111\ : Span4Mux_v
    port map (
            O => \N__32123\,
            I => \N__32117\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__32120\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__32117\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6108\ : CEMux
    port map (
            O => \N__32112\,
            I => \N__32108\
        );

    \I__6107\ : CEMux
    port map (
            O => \N__32111\,
            I => \N__32102\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__32108\,
            I => \N__32097\
        );

    \I__6105\ : CEMux
    port map (
            O => \N__32107\,
            I => \N__32094\
        );

    \I__6104\ : CEMux
    port map (
            O => \N__32106\,
            I => \N__32091\
        );

    \I__6103\ : CEMux
    port map (
            O => \N__32105\,
            I => \N__32088\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32085\
        );

    \I__6101\ : CEMux
    port map (
            O => \N__32101\,
            I => \N__32075\
        );

    \I__6100\ : CEMux
    port map (
            O => \N__32100\,
            I => \N__32072\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__32097\,
            I => \N__32062\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__32062\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32057\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__32088\,
            I => \N__32057\
        );

    \I__6095\ : Span4Mux_h
    port map (
            O => \N__32085\,
            I => \N__32054\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32042\
        );

    \I__6093\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32042\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32042\
        );

    \I__6091\ : CEMux
    port map (
            O => \N__32081\,
            I => \N__32039\
        );

    \I__6090\ : CEMux
    port map (
            O => \N__32080\,
            I => \N__32036\
        );

    \I__6089\ : CEMux
    port map (
            O => \N__32079\,
            I => \N__32033\
        );

    \I__6088\ : CEMux
    port map (
            O => \N__32078\,
            I => \N__32030\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__32075\,
            I => \N__32022\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__32072\,
            I => \N__32019\
        );

    \I__6085\ : CEMux
    port map (
            O => \N__32071\,
            I => \N__32011\
        );

    \I__6084\ : CEMux
    port map (
            O => \N__32070\,
            I => \N__32008\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32001\
        );

    \I__6082\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32001\
        );

    \I__6081\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32001\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__32062\,
            I => \N__31994\
        );

    \I__6079\ : Span4Mux_v
    port map (
            O => \N__32057\,
            I => \N__31994\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__32054\,
            I => \N__31994\
        );

    \I__6077\ : InMux
    port map (
            O => \N__32053\,
            I => \N__31985\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32052\,
            I => \N__31985\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32051\,
            I => \N__31985\
        );

    \I__6074\ : InMux
    port map (
            O => \N__32050\,
            I => \N__31985\
        );

    \I__6073\ : CEMux
    port map (
            O => \N__32049\,
            I => \N__31981\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__31978\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__32039\,
            I => \N__31975\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__31968\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__32033\,
            I => \N__31968\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__32030\,
            I => \N__31968\
        );

    \I__6067\ : CEMux
    port map (
            O => \N__32029\,
            I => \N__31953\
        );

    \I__6066\ : InMux
    port map (
            O => \N__32028\,
            I => \N__31944\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32027\,
            I => \N__31944\
        );

    \I__6064\ : InMux
    port map (
            O => \N__32026\,
            I => \N__31944\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32025\,
            I => \N__31944\
        );

    \I__6062\ : Span4Mux_v
    port map (
            O => \N__32022\,
            I => \N__31939\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__32019\,
            I => \N__31939\
        );

    \I__6060\ : CEMux
    port map (
            O => \N__32018\,
            I => \N__31936\
        );

    \I__6059\ : InMux
    port map (
            O => \N__32017\,
            I => \N__31927\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31927\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31927\
        );

    \I__6056\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31927\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__32011\,
            I => \N__31924\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__32008\,
            I => \N__31921\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31918\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__31994\,
            I => \N__31913\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__31985\,
            I => \N__31913\
        );

    \I__6050\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31910\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__31981\,
            I => \N__31907\
        );

    \I__6048\ : Span4Mux_h
    port map (
            O => \N__31978\,
            I => \N__31902\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__31975\,
            I => \N__31902\
        );

    \I__6046\ : Span4Mux_v
    port map (
            O => \N__31968\,
            I => \N__31899\
        );

    \I__6045\ : InMux
    port map (
            O => \N__31967\,
            I => \N__31890\
        );

    \I__6044\ : InMux
    port map (
            O => \N__31966\,
            I => \N__31890\
        );

    \I__6043\ : InMux
    port map (
            O => \N__31965\,
            I => \N__31890\
        );

    \I__6042\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31890\
        );

    \I__6041\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31881\
        );

    \I__6040\ : InMux
    port map (
            O => \N__31962\,
            I => \N__31881\
        );

    \I__6039\ : InMux
    port map (
            O => \N__31961\,
            I => \N__31881\
        );

    \I__6038\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31881\
        );

    \I__6037\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31872\
        );

    \I__6036\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31872\
        );

    \I__6035\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31872\
        );

    \I__6034\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31872\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__31953\,
            I => \N__31865\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31865\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__31939\,
            I => \N__31865\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__31936\,
            I => \N__31856\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__31927\,
            I => \N__31856\
        );

    \I__6028\ : Span4Mux_v
    port map (
            O => \N__31924\,
            I => \N__31856\
        );

    \I__6027\ : Span4Mux_v
    port map (
            O => \N__31921\,
            I => \N__31856\
        );

    \I__6026\ : Span4Mux_h
    port map (
            O => \N__31918\,
            I => \N__31851\
        );

    \I__6025\ : Span4Mux_h
    port map (
            O => \N__31913\,
            I => \N__31851\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__31910\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6023\ : Odrv12
    port map (
            O => \N__31907\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6022\ : Odrv4
    port map (
            O => \N__31902\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__31899\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__31890\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__31881\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6018\ : LocalMux
    port map (
            O => \N__31872\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6017\ : Odrv4
    port map (
            O => \N__31865\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__31856\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6015\ : Odrv4
    port map (
            O => \N__31851\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__6014\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31827\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__31827\,
            I => \N__31823\
        );

    \I__6012\ : InMux
    port map (
            O => \N__31826\,
            I => \N__31819\
        );

    \I__6011\ : Span4Mux_h
    port map (
            O => \N__31823\,
            I => \N__31816\
        );

    \I__6010\ : InMux
    port map (
            O => \N__31822\,
            I => \N__31813\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__31819\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__31816\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__31813\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6006\ : InMux
    port map (
            O => \N__31806\,
            I => \N__31803\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__31803\,
            I => \N__31800\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__31800\,
            I => \phase_controller_inst2.start_timer_hc_0_sqmuxa\
        );

    \I__6003\ : IoInMux
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__6001\ : Span4Mux_s2_v
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__31788\,
            I => \N__31785\
        );

    \I__5999\ : Span4Mux_v
    port map (
            O => \N__31785\,
            I => \N__31780\
        );

    \I__5998\ : InMux
    port map (
            O => \N__31784\,
            I => \N__31775\
        );

    \I__5997\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31775\
        );

    \I__5996\ : Odrv4
    port map (
            O => \N__31780\,
            I => s1_phy_c
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__31775\,
            I => s1_phy_c
        );

    \I__5994\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31761\
        );

    \I__5993\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31761\
        );

    \I__5992\ : InMux
    port map (
            O => \N__31768\,
            I => \N__31761\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__31761\,
            I => \N__31756\
        );

    \I__5990\ : InMux
    port map (
            O => \N__31760\,
            I => \N__31752\
        );

    \I__5989\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31749\
        );

    \I__5988\ : Span4Mux_v
    port map (
            O => \N__31756\,
            I => \N__31746\
        );

    \I__5987\ : InMux
    port map (
            O => \N__31755\,
            I => \N__31743\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__31752\,
            I => state_3
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__31749\,
            I => state_3
        );

    \I__5984\ : Odrv4
    port map (
            O => \N__31746\,
            I => state_3
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__31743\,
            I => state_3
        );

    \I__5982\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__31731\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__5979\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31722\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__31722\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__5977\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31716\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__31716\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__5975\ : CascadeMux
    port map (
            O => \N__31713\,
            I => \N__31710\
        );

    \I__5974\ : InMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__31707\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__31704\,
            I => \N__31701\
        );

    \I__5971\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31698\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__31698\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__5969\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__5968\ : LocalMux
    port map (
            O => \N__31692\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__31689\,
            I => \N__31686\
        );

    \I__5966\ : InMux
    port map (
            O => \N__31686\,
            I => \N__31683\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__31683\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__5964\ : InMux
    port map (
            O => \N__31680\,
            I => \N__31677\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__31674\,
            I => \N__31671\
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__31671\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__5960\ : InMux
    port map (
            O => \N__31668\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__5959\ : CascadeMux
    port map (
            O => \N__31665\,
            I => \N__31662\
        );

    \I__5958\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31659\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__31659\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__5956\ : InMux
    port map (
            O => \N__31656\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__5955\ : InMux
    port map (
            O => \N__31653\,
            I => \N__31650\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__5953\ : Span4Mux_h
    port map (
            O => \N__31647\,
            I => \N__31644\
        );

    \I__5952\ : Odrv4
    port map (
            O => \N__31644\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__5951\ : InMux
    port map (
            O => \N__31641\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__5950\ : InMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__31635\,
            I => \N__31632\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__31632\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__5947\ : InMux
    port map (
            O => \N__31629\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__5946\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31623\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__31620\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__5943\ : InMux
    port map (
            O => \N__31617\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__5942\ : InMux
    port map (
            O => \N__31614\,
            I => \N__31611\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__31611\,
            I => \N__31608\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__31608\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__5939\ : InMux
    port map (
            O => \N__31605\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__5938\ : InMux
    port map (
            O => \N__31602\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__5937\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31596\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__31596\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__5935\ : InMux
    port map (
            O => \N__31593\,
            I => \N__31590\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__31590\,
            I => \N__31587\
        );

    \I__5933\ : Span4Mux_v
    port map (
            O => \N__31587\,
            I => \N__31584\
        );

    \I__5932\ : Odrv4
    port map (
            O => \N__31584\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__5931\ : InMux
    port map (
            O => \N__31581\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__5930\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31575\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__31575\,
            I => \N__31572\
        );

    \I__5928\ : Span4Mux_v
    port map (
            O => \N__31572\,
            I => \N__31569\
        );

    \I__5927\ : Odrv4
    port map (
            O => \N__31569\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__5926\ : InMux
    port map (
            O => \N__31566\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__5925\ : InMux
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__31557\,
            I => \N__31554\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__31554\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__5921\ : InMux
    port map (
            O => \N__31551\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__5920\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__5918\ : Span4Mux_h
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__31539\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__5916\ : InMux
    port map (
            O => \N__31536\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__5915\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__31530\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__5913\ : InMux
    port map (
            O => \N__31527\,
            I => \bfn_12_20_0_\
        );

    \I__5912\ : CascadeMux
    port map (
            O => \N__31524\,
            I => \N__31521\
        );

    \I__5911\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31518\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__31518\,
            I => \N__31515\
        );

    \I__5909\ : Odrv12
    port map (
            O => \N__31515\,
            I => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__31512\,
            I => \N__31509\
        );

    \I__5907\ : InMux
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__31506\,
            I => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\
        );

    \I__5905\ : CascadeMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__5904\ : InMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__31497\,
            I => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\
        );

    \I__5902\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31484\
        );

    \I__5901\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31484\
        );

    \I__5900\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31484\
        );

    \I__5899\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31481\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__31484\,
            I => \N__31478\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__31481\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__31478\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31473\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__5894\ : InMux
    port map (
            O => \N__31470\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__31467\,
            I => \N__31463\
        );

    \I__5892\ : CascadeMux
    port map (
            O => \N__31466\,
            I => \N__31459\
        );

    \I__5891\ : InMux
    port map (
            O => \N__31463\,
            I => \N__31452\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31452\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31452\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N__31448\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31445\
        );

    \I__5886\ : Span4Mux_h
    port map (
            O => \N__31448\,
            I => \N__31442\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__31445\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__31442\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__5883\ : CascadeMux
    port map (
            O => \N__31437\,
            I => \N__31433\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31429\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31426\
        );

    \I__5880\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31423\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__31429\,
            I => \il_max_comp1_D2\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__31426\,
            I => \il_max_comp1_D2\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31423\,
            I => \il_max_comp1_D2\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__31416\,
            I => \N__31413\
        );

    \I__5875\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31407\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__31407\,
            I => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\
        );

    \I__5872\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31401\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__5870\ : Odrv4
    port map (
            O => \N__31398\,
            I => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__31395\,
            I => \N__31392\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31389\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31389\,
            I => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\
        );

    \I__5866\ : CascadeMux
    port map (
            O => \N__31386\,
            I => \N__31383\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31380\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31377\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__31377\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__31374\,
            I => \N__31371\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31365\
        );

    \I__5860\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31365\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31361\
        );

    \I__5858\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31358\
        );

    \I__5857\ : Span4Mux_h
    port map (
            O => \N__31361\,
            I => \N__31355\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__31358\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__5855\ : Odrv4
    port map (
            O => \N__31355\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__5854\ : InMux
    port map (
            O => \N__31350\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__5853\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31341\
        );

    \I__5852\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31341\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__31341\,
            I => \N__31337\
        );

    \I__5850\ : InMux
    port map (
            O => \N__31340\,
            I => \N__31334\
        );

    \I__5849\ : Span4Mux_h
    port map (
            O => \N__31337\,
            I => \N__31331\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__31334\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__5847\ : Odrv4
    port map (
            O => \N__31331\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__5846\ : InMux
    port map (
            O => \N__31326\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__5845\ : CascadeMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__5844\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31314\
        );

    \I__5843\ : InMux
    port map (
            O => \N__31319\,
            I => \N__31314\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__31314\,
            I => \N__31310\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31307\
        );

    \I__5840\ : Span4Mux_h
    port map (
            O => \N__31310\,
            I => \N__31304\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__31307\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__5838\ : Odrv4
    port map (
            O => \N__31304\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__5837\ : InMux
    port map (
            O => \N__31299\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__5836\ : InMux
    port map (
            O => \N__31296\,
            I => \N__31289\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31295\,
            I => \N__31289\
        );

    \I__5834\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31286\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__31289\,
            I => \N__31283\
        );

    \I__5832\ : LocalMux
    port map (
            O => \N__31286\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__5831\ : Odrv4
    port map (
            O => \N__31283\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__5830\ : InMux
    port map (
            O => \N__31278\,
            I => \bfn_12_13_0_\
        );

    \I__5829\ : InMux
    port map (
            O => \N__31275\,
            I => \N__31271\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__31274\,
            I => \N__31268\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__31271\,
            I => \N__31264\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31268\,
            I => \N__31261\
        );

    \I__5825\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31258\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__31264\,
            I => \N__31253\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31261\,
            I => \N__31253\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31258\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__31253\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31248\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__31245\,
            I => \N__31242\
        );

    \I__5818\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31238\
        );

    \I__5817\ : InMux
    port map (
            O => \N__31241\,
            I => \N__31234\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__31238\,
            I => \N__31231\
        );

    \I__5815\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31228\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31234\,
            I => \N__31225\
        );

    \I__5813\ : Span4Mux_h
    port map (
            O => \N__31231\,
            I => \N__31222\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__31228\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__5811\ : Odrv4
    port map (
            O => \N__31225\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__31222\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31215\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31209\,
            I => \N__31203\
        );

    \I__5806\ : InMux
    port map (
            O => \N__31208\,
            I => \N__31203\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__31203\,
            I => \N__31199\
        );

    \I__5804\ : InMux
    port map (
            O => \N__31202\,
            I => \N__31196\
        );

    \I__5803\ : Span4Mux_h
    port map (
            O => \N__31199\,
            I => \N__31193\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__31196\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__31193\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__5800\ : InMux
    port map (
            O => \N__31188\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__5799\ : InMux
    port map (
            O => \N__31185\,
            I => \N__31179\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31179\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__31179\,
            I => \N__31175\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31172\
        );

    \I__5795\ : Span4Mux_h
    port map (
            O => \N__31175\,
            I => \N__31169\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31172\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5793\ : Odrv4
    port map (
            O => \N__31169\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31164\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31157\
        );

    \I__5790\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31154\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31157\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__31154\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31149\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__5786\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31142\
        );

    \I__5785\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31139\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__31142\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__31139\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31134\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31127\
        );

    \I__5780\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31124\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31127\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__31124\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31119\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__31116\,
            I => \N__31113\
        );

    \I__5775\ : InMux
    port map (
            O => \N__31113\,
            I => \N__31107\
        );

    \I__5774\ : InMux
    port map (
            O => \N__31112\,
            I => \N__31107\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__31107\,
            I => \N__31103\
        );

    \I__5772\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31100\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__31103\,
            I => \N__31097\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31100\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__31097\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31092\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__5767\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31082\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31082\
        );

    \I__5765\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31079\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__31082\,
            I => \N__31076\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__31079\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5762\ : Odrv12
    port map (
            O => \N__31076\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__5761\ : InMux
    port map (
            O => \N__31071\,
            I => \bfn_12_12_0_\
        );

    \I__5760\ : InMux
    port map (
            O => \N__31068\,
            I => \N__31062\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31067\,
            I => \N__31062\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__31062\,
            I => \N__31058\
        );

    \I__5757\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31055\
        );

    \I__5756\ : Span4Mux_h
    port map (
            O => \N__31058\,
            I => \N__31052\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__31055\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__31052\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__5753\ : InMux
    port map (
            O => \N__31047\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__31044\,
            I => \N__31041\
        );

    \I__5751\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31035\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31040\,
            I => \N__31035\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__31035\,
            I => \N__31031\
        );

    \I__5748\ : InMux
    port map (
            O => \N__31034\,
            I => \N__31028\
        );

    \I__5747\ : Span4Mux_v
    port map (
            O => \N__31031\,
            I => \N__31025\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__31028\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__31025\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__5744\ : InMux
    port map (
            O => \N__31020\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__5743\ : InMux
    port map (
            O => \N__31017\,
            I => \N__31011\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31016\,
            I => \N__31011\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__31011\,
            I => \N__31007\
        );

    \I__5740\ : InMux
    port map (
            O => \N__31010\,
            I => \N__31004\
        );

    \I__5739\ : Span4Mux_h
    port map (
            O => \N__31007\,
            I => \N__31001\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__31004\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__5737\ : Odrv4
    port map (
            O => \N__31001\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__5736\ : InMux
    port map (
            O => \N__30996\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__30993\,
            I => \N__30990\
        );

    \I__5734\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30984\
        );

    \I__5733\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30984\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__30984\,
            I => \N__30980\
        );

    \I__5731\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30977\
        );

    \I__5730\ : Span4Mux_v
    port map (
            O => \N__30980\,
            I => \N__30974\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__30977\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__5728\ : Odrv4
    port map (
            O => \N__30974\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__5727\ : InMux
    port map (
            O => \N__30969\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__5726\ : InMux
    port map (
            O => \N__30966\,
            I => \N__30962\
        );

    \I__5725\ : InMux
    port map (
            O => \N__30965\,
            I => \N__30959\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__30962\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__30959\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5722\ : InMux
    port map (
            O => \N__30954\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__5721\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30947\
        );

    \I__5720\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30944\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__30947\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__30944\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5717\ : InMux
    port map (
            O => \N__30939\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__5716\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30932\
        );

    \I__5715\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30929\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__30932\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__30929\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5712\ : InMux
    port map (
            O => \N__30924\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__5711\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30917\
        );

    \I__5710\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30914\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__30917\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5708\ : LocalMux
    port map (
            O => \N__30914\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5707\ : InMux
    port map (
            O => \N__30909\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__5706\ : InMux
    port map (
            O => \N__30906\,
            I => \N__30902\
        );

    \I__5705\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30899\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__30902\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__30899\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5702\ : InMux
    port map (
            O => \N__30894\,
            I => \bfn_12_11_0_\
        );

    \I__5701\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30887\
        );

    \I__5700\ : InMux
    port map (
            O => \N__30890\,
            I => \N__30884\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__30887\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__30884\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5697\ : InMux
    port map (
            O => \N__30879\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__5696\ : InMux
    port map (
            O => \N__30876\,
            I => \N__30872\
        );

    \I__5695\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30869\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__30872\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__30869\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5692\ : InMux
    port map (
            O => \N__30864\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__5691\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30857\
        );

    \I__5690\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30854\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__30857\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__30854\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5687\ : InMux
    port map (
            O => \N__30849\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__5686\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30843\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__30843\,
            I => \N__30840\
        );

    \I__5684\ : Span4Mux_h
    port map (
            O => \N__30840\,
            I => \N__30837\
        );

    \I__5683\ : Odrv4
    port map (
            O => \N__30837\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__30834\,
            I => \N__30831\
        );

    \I__5681\ : InMux
    port map (
            O => \N__30831\,
            I => \N__30828\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30825\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__30825\,
            I => \N__30822\
        );

    \I__5678\ : Odrv4
    port map (
            O => \N__30822\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__5677\ : InMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__5675\ : Span4Mux_h
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__30810\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__5673\ : CascadeMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__5672\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__30801\,
            I => \N__30798\
        );

    \I__5670\ : Span4Mux_v
    port map (
            O => \N__30798\,
            I => \N__30795\
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__30795\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__5668\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30789\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__30789\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__5666\ : CascadeMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__5665\ : InMux
    port map (
            O => \N__30783\,
            I => \N__30779\
        );

    \I__5664\ : InMux
    port map (
            O => \N__30782\,
            I => \N__30776\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__30779\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__30776\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__5661\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30768\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__30768\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__5659\ : InMux
    port map (
            O => \N__30765\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_28\
        );

    \I__5658\ : InMux
    port map (
            O => \N__30762\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__5657\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30753\
        );

    \I__5656\ : InMux
    port map (
            O => \N__30758\,
            I => \N__30753\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__30753\,
            I => \N__30750\
        );

    \I__5654\ : Odrv12
    port map (
            O => \N__30750\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__5653\ : InMux
    port map (
            O => \N__30747\,
            I => \N__30744\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__30744\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__30741\,
            I => \N__30737\
        );

    \I__5650\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30733\
        );

    \I__5649\ : InMux
    port map (
            O => \N__30737\,
            I => \N__30730\
        );

    \I__5648\ : InMux
    port map (
            O => \N__30736\,
            I => \N__30727\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__30733\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__30730\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__30727\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__5644\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30716\
        );

    \I__5643\ : InMux
    port map (
            O => \N__30719\,
            I => \N__30713\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__30716\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__30713\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5640\ : InMux
    port map (
            O => \N__30708\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__5639\ : CascadeMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__5638\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__30699\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\
        );

    \I__5636\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30692\
        );

    \I__5635\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30689\
        );

    \I__5634\ : LocalMux
    port map (
            O => \N__30692\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__30689\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5632\ : InMux
    port map (
            O => \N__30684\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__5631\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30677\
        );

    \I__5630\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30674\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__30677\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__30674\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5627\ : InMux
    port map (
            O => \N__30669\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__5626\ : InMux
    port map (
            O => \N__30666\,
            I => \N__30662\
        );

    \I__5625\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30659\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30656\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__30659\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5622\ : Odrv4
    port map (
            O => \N__30656\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__5621\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30648\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__30648\,
            I => \N__30645\
        );

    \I__5619\ : Span4Mux_h
    port map (
            O => \N__30645\,
            I => \N__30642\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__30639\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__5616\ : CascadeMux
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__5615\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30630\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__30627\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__5612\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30621\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__30621\,
            I => \N__30617\
        );

    \I__5610\ : InMux
    port map (
            O => \N__30620\,
            I => \N__30614\
        );

    \I__5609\ : Span4Mux_v
    port map (
            O => \N__30617\,
            I => \N__30611\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__30614\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__30611\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__30606\,
            I => \N__30603\
        );

    \I__5605\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30600\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__30600\,
            I => \N__30597\
        );

    \I__5603\ : Odrv12
    port map (
            O => \N__30597\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__5602\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30591\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__30591\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__5600\ : InMux
    port map (
            O => \N__30588\,
            I => \N__30585\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__30585\,
            I => \N__30582\
        );

    \I__5598\ : Odrv12
    port map (
            O => \N__30582\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__5597\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30575\
        );

    \I__5596\ : InMux
    port map (
            O => \N__30578\,
            I => \N__30572\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__30575\,
            I => \N__30569\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__30572\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__30569\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__30564\,
            I => \N__30561\
        );

    \I__5591\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30558\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__30558\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__5589\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30552\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__5587\ : Odrv4
    port map (
            O => \N__30549\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__5586\ : CascadeMux
    port map (
            O => \N__30546\,
            I => \N__30543\
        );

    \I__5585\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__30540\,
            I => \N__30537\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__5582\ : Odrv4
    port map (
            O => \N__30534\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__5581\ : InMux
    port map (
            O => \N__30531\,
            I => \N__30528\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__30525\,
            I => \N__30522\
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__30522\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__5576\ : InMux
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__30513\,
            I => \N__30510\
        );

    \I__5574\ : Span4Mux_v
    port map (
            O => \N__30510\,
            I => \N__30507\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__30507\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__5572\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30501\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__30501\,
            I => \N__30498\
        );

    \I__5570\ : Odrv4
    port map (
            O => \N__30498\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__5568\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30489\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__30486\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__5565\ : InMux
    port map (
            O => \N__30483\,
            I => \N__30480\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__30480\,
            I => \N__30477\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__30477\,
            I => \N__30474\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__30474\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__5560\ : InMux
    port map (
            O => \N__30468\,
            I => \N__30465\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__30465\,
            I => \N__30462\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__5557\ : Odrv4
    port map (
            O => \N__30459\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__5556\ : InMux
    port map (
            O => \N__30456\,
            I => \N__30453\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5554\ : Span4Mux_v
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__5553\ : Odrv4
    port map (
            O => \N__30447\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__5552\ : CascadeMux
    port map (
            O => \N__30444\,
            I => \N__30441\
        );

    \I__5551\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30435\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__30435\,
            I => \N__30432\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__30432\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30425\
        );

    \I__5546\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30422\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__30425\,
            I => \N__30419\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__30422\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5543\ : Odrv4
    port map (
            O => \N__30419\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__30408\,
            I => \N__30405\
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__30405\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__5537\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30396\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__5535\ : Odrv4
    port map (
            O => \N__30393\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__5534\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30387\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30384\
        );

    \I__5532\ : Odrv12
    port map (
            O => \N__30384\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30377\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30374\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30371\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__30374\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5527\ : Odrv4
    port map (
            O => \N__30371\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__5525\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30360\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__5523\ : InMux
    port map (
            O => \N__30357\,
            I => \N__30353\
        );

    \I__5522\ : InMux
    port map (
            O => \N__30356\,
            I => \N__30350\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__30353\,
            I => \N__30347\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__30350\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5519\ : Odrv4
    port map (
            O => \N__30347\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__5518\ : InMux
    port map (
            O => \N__30342\,
            I => \N__30339\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__5516\ : Span4Mux_v
    port map (
            O => \N__30336\,
            I => \N__30333\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__30333\,
            I => \N__30330\
        );

    \I__5514\ : Span4Mux_h
    port map (
            O => \N__30330\,
            I => \N__30327\
        );

    \I__5513\ : Odrv4
    port map (
            O => \N__30327\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__5512\ : CascadeMux
    port map (
            O => \N__30324\,
            I => \N__30321\
        );

    \I__5511\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__30315\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__5508\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30309\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__5506\ : Span4Mux_h
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__5505\ : Odrv4
    port map (
            O => \N__30303\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30297\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30297\,
            I => \N__30293\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30290\
        );

    \I__5501\ : Span4Mux_v
    port map (
            O => \N__30293\,
            I => \N__30287\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__30290\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__30287\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__5498\ : CascadeMux
    port map (
            O => \N__30282\,
            I => \N__30279\
        );

    \I__5497\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30276\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__30276\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__5495\ : InMux
    port map (
            O => \N__30273\,
            I => \N__30270\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__30267\,
            I => \N__30264\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__30264\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__5491\ : InMux
    port map (
            O => \N__30261\,
            I => \N__30257\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30254\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30251\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__30254\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5487\ : Odrv4
    port map (
            O => \N__30251\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__5486\ : CascadeMux
    port map (
            O => \N__30246\,
            I => \N__30243\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30240\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__30240\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__5483\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30234\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__30234\,
            I => \N__30231\
        );

    \I__5481\ : Span4Mux_h
    port map (
            O => \N__30231\,
            I => \N__30228\
        );

    \I__5480\ : Odrv4
    port map (
            O => \N__30228\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__5479\ : InMux
    port map (
            O => \N__30225\,
            I => \N__30222\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30222\,
            I => \N__30218\
        );

    \I__5477\ : InMux
    port map (
            O => \N__30221\,
            I => \N__30215\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__30218\,
            I => \N__30212\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30215\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5474\ : Odrv4
    port map (
            O => \N__30212\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__5473\ : CascadeMux
    port map (
            O => \N__30207\,
            I => \N__30204\
        );

    \I__5472\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30201\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30201\,
            I => \N__30198\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__30198\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__5467\ : Odrv12
    port map (
            O => \N__30189\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__5466\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30182\
        );

    \I__5465\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30179\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30176\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__30179\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__30176\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__5461\ : CascadeMux
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__5460\ : InMux
    port map (
            O => \N__30168\,
            I => \N__30165\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30165\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__30162\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\
        );

    \I__5457\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__30156\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30141\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30152\,
            I => \N__30141\
        );

    \I__5453\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30141\
        );

    \I__5452\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30141\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__30141\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__30138\,
            I => \N__30133\
        );

    \I__5449\ : CascadeMux
    port map (
            O => \N__30137\,
            I => \N__30130\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30136\,
            I => \N__30125\
        );

    \I__5447\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30116\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30130\,
            I => \N__30116\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30129\,
            I => \N__30116\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30116\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__30125\,
            I => \N__30113\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__30116\,
            I => \N__30108\
        );

    \I__5441\ : Span4Mux_v
    port map (
            O => \N__30113\,
            I => \N__30108\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__30108\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30102\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30102\,
            I => \N__30099\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__30099\,
            I => \N__30096\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__30096\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__30093\,
            I => \N__30090\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30087\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30087\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30084\,
            I => \N__30081\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30081\,
            I => \N__30078\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__30078\,
            I => \N__30075\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__30075\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__5428\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30068\
        );

    \I__5427\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30065\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__30068\,
            I => \N__30062\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__30065\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5424\ : Odrv4
    port map (
            O => \N__30062\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__30057\,
            I => \N__30054\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30051\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__30051\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30048\,
            I => \N__30045\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30045\,
            I => \N__30042\
        );

    \I__5418\ : Span4Mux_h
    port map (
            O => \N__30042\,
            I => \N__30039\
        );

    \I__5417\ : Odrv4
    port map (
            O => \N__30039\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30032\
        );

    \I__5415\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30029\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30026\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30023\
        );

    \I__5412\ : Span4Mux_v
    port map (
            O => \N__30026\,
            I => \N__30020\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__30023\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__30020\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__5409\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__5408\ : InMux
    port map (
            O => \N__30012\,
            I => \N__30009\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__30009\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30006\,
            I => \N__30003\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__30003\,
            I => \N__30000\
        );

    \I__5404\ : Span4Mux_v
    port map (
            O => \N__30000\,
            I => \N__29997\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__29997\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__5402\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29990\
        );

    \I__5401\ : InMux
    port map (
            O => \N__29993\,
            I => \N__29987\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29984\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__29987\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__29984\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__29979\,
            I => \N__29976\
        );

    \I__5396\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__29973\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__5394\ : InMux
    port map (
            O => \N__29970\,
            I => \N__29966\
        );

    \I__5393\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29963\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__29966\,
            I => \N__29960\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__29963\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__29960\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__5389\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29952\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29949\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__29949\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__29946\,
            I => \N__29943\
        );

    \I__5385\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29940\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__29940\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__5383\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29933\
        );

    \I__5382\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29929\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__29933\,
            I => \N__29926\
        );

    \I__5380\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29923\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__29929\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__5378\ : Odrv4
    port map (
            O => \N__29926\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__29923\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__29916\,
            I => \N__29913\
        );

    \I__5375\ : InMux
    port map (
            O => \N__29913\,
            I => \N__29910\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__29910\,
            I => \N__29907\
        );

    \I__5373\ : Span4Mux_h
    port map (
            O => \N__29907\,
            I => \N__29903\
        );

    \I__5372\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29900\
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__29903\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__29900\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__5369\ : InMux
    port map (
            O => \N__29895\,
            I => \N__29892\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__5367\ : Odrv12
    port map (
            O => \N__29889\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__29886\,
            I => \N__29882\
        );

    \I__5365\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29877\
        );

    \I__5364\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29874\
        );

    \I__5363\ : CascadeMux
    port map (
            O => \N__29881\,
            I => \N__29869\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__29880\,
            I => \N__29863\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29858\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__29874\,
            I => \N__29858\
        );

    \I__5359\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29855\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__29872\,
            I => \N__29852\
        );

    \I__5357\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29843\
        );

    \I__5356\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29843\
        );

    \I__5355\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29843\
        );

    \I__5354\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29843\
        );

    \I__5353\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29840\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__29858\,
            I => \N__29835\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29835\
        );

    \I__5350\ : InMux
    port map (
            O => \N__29852\,
            I => \N__29832\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__29843\,
            I => \N__29824\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__29840\,
            I => \N__29824\
        );

    \I__5347\ : Span4Mux_v
    port map (
            O => \N__29835\,
            I => \N__29821\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29818\
        );

    \I__5345\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29815\
        );

    \I__5344\ : InMux
    port map (
            O => \N__29830\,
            I => \N__29810\
        );

    \I__5343\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29810\
        );

    \I__5342\ : Span4Mux_v
    port map (
            O => \N__29824\,
            I => \N__29807\
        );

    \I__5341\ : Span4Mux_s2_v
    port map (
            O => \N__29821\,
            I => \N__29804\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__29818\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__29815\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__29810\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5337\ : Odrv4
    port map (
            O => \N__29807\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__29804\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__5335\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__29790\,
            I => \N__29787\
        );

    \I__5333\ : Odrv12
    port map (
            O => \N__29787\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__5332\ : CascadeMux
    port map (
            O => \N__29784\,
            I => \N__29781\
        );

    \I__5331\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29777\
        );

    \I__5330\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29773\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__29777\,
            I => \N__29770\
        );

    \I__5328\ : InMux
    port map (
            O => \N__29776\,
            I => \N__29767\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__29773\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__5326\ : Odrv4
    port map (
            O => \N__29770\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__29767\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__5324\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29757\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__29757\,
            I => \N__29754\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__29754\,
            I => \N__29750\
        );

    \I__5321\ : InMux
    port map (
            O => \N__29753\,
            I => \N__29747\
        );

    \I__5320\ : Odrv4
    port map (
            O => \N__29750\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__29747\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__5318\ : InMux
    port map (
            O => \N__29742\,
            I => \N__29739\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__29739\,
            I => \N__29736\
        );

    \I__5316\ : Odrv12
    port map (
            O => \N__29736\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__5315\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29729\
        );

    \I__5314\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29726\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__29729\,
            I => \N__29723\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29720\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__29723\,
            I => \N__29715\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__29720\,
            I => \N__29715\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__29715\,
            I => \N__29710\
        );

    \I__5308\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29707\
        );

    \I__5307\ : InMux
    port map (
            O => \N__29713\,
            I => \N__29704\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__29710\,
            I => \N__29701\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__29707\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__29704\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5303\ : Odrv4
    port map (
            O => \N__29701\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5302\ : ClkMux
    port map (
            O => \N__29694\,
            I => \N__29688\
        );

    \I__5301\ : ClkMux
    port map (
            O => \N__29693\,
            I => \N__29688\
        );

    \I__5300\ : GlobalMux
    port map (
            O => \N__29688\,
            I => \N__29685\
        );

    \I__5299\ : gio2CtrlBuf
    port map (
            O => \N__29685\,
            I => delay_hc_input_c_g
        );

    \I__5298\ : InMux
    port map (
            O => \N__29682\,
            I => \N__29677\
        );

    \I__5297\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29673\
        );

    \I__5296\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29670\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__29677\,
            I => \N__29667\
        );

    \I__5294\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29664\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__29673\,
            I => \N__29661\
        );

    \I__5292\ : InMux
    port map (
            O => \N__29670\,
            I => \N__29658\
        );

    \I__5291\ : Span4Mux_v
    port map (
            O => \N__29667\,
            I => \N__29655\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__29664\,
            I => \N__29648\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__29661\,
            I => \N__29648\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__29658\,
            I => \N__29648\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__29655\,
            I => \N__29645\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__29648\,
            I => \N__29642\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__29645\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__29642\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__5283\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29632\
        );

    \I__5282\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29629\
        );

    \I__5281\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29626\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__29632\,
            I => \N__29623\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__29629\,
            I => \N__29620\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__29626\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__5277\ : Odrv12
    port map (
            O => \N__29623\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__29620\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__5275\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__29610\,
            I => \N__29607\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__29607\,
            I => \N__29604\
        );

    \I__5272\ : Span4Mux_v
    port map (
            O => \N__29604\,
            I => \N__29601\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__29601\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__5270\ : CascadeMux
    port map (
            O => \N__29598\,
            I => \N__29595\
        );

    \I__5269\ : InMux
    port map (
            O => \N__29595\,
            I => \N__29592\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__29592\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__5267\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29583\
        );

    \I__5266\ : InMux
    port map (
            O => \N__29588\,
            I => \N__29583\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__29583\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__5264\ : InMux
    port map (
            O => \N__29580\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__5263\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29574\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__29574\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__5261\ : InMux
    port map (
            O => \N__29571\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__5260\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__29565\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__5258\ : InMux
    port map (
            O => \N__29562\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__5257\ : InMux
    port map (
            O => \N__29559\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__5256\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__29553\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__5254\ : InMux
    port map (
            O => \N__29550\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__5253\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__29544\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__5251\ : InMux
    port map (
            O => \N__29541\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__5250\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__29535\,
            I => \N__29532\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__29532\,
            I => \N__29529\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__29529\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__5246\ : InMux
    port map (
            O => \N__29526\,
            I => \bfn_11_25_0_\
        );

    \I__5245\ : InMux
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__29520\,
            I => \N__29517\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__29517\,
            I => \N__29514\
        );

    \I__5242\ : Odrv4
    port map (
            O => \N__29514\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__5241\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__5238\ : Odrv4
    port map (
            O => \N__29502\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__5237\ : InMux
    port map (
            O => \N__29499\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__5236\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29493\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__5234\ : Odrv12
    port map (
            O => \N__29490\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__5231\ : Odrv12
    port map (
            O => \N__29481\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__5230\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29475\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__29475\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__5228\ : InMux
    port map (
            O => \N__29472\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__5227\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29466\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__29466\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__5225\ : InMux
    port map (
            O => \N__29463\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__5224\ : InMux
    port map (
            O => \N__29460\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__5223\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29451\
        );

    \I__5221\ : Span12Mux_v
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__5220\ : Odrv12
    port map (
            O => \N__29448\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__5219\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__29442\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__29436\,
            I => \N__29433\
        );

    \I__5215\ : Span4Mux_v
    port map (
            O => \N__29433\,
            I => \N__29430\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__29430\,
            I => \N__29427\
        );

    \I__5213\ : Odrv4
    port map (
            O => \N__29427\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29424\,
            I => \N__29421\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__29421\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__5210\ : InMux
    port map (
            O => \N__29418\,
            I => \N__29415\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__29409\,
            I => \N__29406\
        );

    \I__5206\ : Odrv4
    port map (
            O => \N__29406\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__5205\ : IoInMux
    port map (
            O => \N__29403\,
            I => \N__29400\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29400\,
            I => \N__29397\
        );

    \I__5203\ : Span4Mux_s3_v
    port map (
            O => \N__29397\,
            I => \N__29394\
        );

    \I__5202\ : Span4Mux_v
    port map (
            O => \N__29394\,
            I => \N__29391\
        );

    \I__5201\ : Odrv4
    port map (
            O => \N__29391\,
            I => s3_phy_c
        );

    \I__5200\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29385\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__29385\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29379\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__29379\,
            I => \N__29376\
        );

    \I__5196\ : Span4Mux_h
    port map (
            O => \N__29376\,
            I => \N__29373\
        );

    \I__5195\ : Odrv4
    port map (
            O => \N__29373\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29370\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__5193\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29364\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__29364\,
            I => \N__29361\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__29361\,
            I => \N__29358\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__29358\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__5189\ : InMux
    port map (
            O => \N__29355\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29352\,
            I => \N__29349\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__29346\,
            I => \N__29343\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__29343\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29340\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__5183\ : InMux
    port map (
            O => \N__29337\,
            I => \N__29334\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__5180\ : Odrv4
    port map (
            O => \N__29328\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29325\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__5178\ : InMux
    port map (
            O => \N__29322\,
            I => \bfn_11_20_0_\
        );

    \I__5177\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29316\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__5175\ : Span4Mux_h
    port map (
            O => \N__29313\,
            I => \N__29310\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__29310\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__5173\ : InMux
    port map (
            O => \N__29307\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29304\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__29298\,
            I => \N__29295\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__29295\,
            I => \N__29292\
        );

    \I__5168\ : Odrv4
    port map (
            O => \N__29292\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29289\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29283\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__29283\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29280\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29271\
        );

    \I__5161\ : LocalMux
    port map (
            O => \N__29271\,
            I => \N__29268\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__29268\,
            I => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29265\,
            I => \N__29262\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29259\
        );

    \I__5157\ : Odrv4
    port map (
            O => \N__29259\,
            I => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\
        );

    \I__5156\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__5154\ : Span4Mux_v
    port map (
            O => \N__29250\,
            I => \N__29247\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__29247\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29244\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__5151\ : CascadeMux
    port map (
            O => \N__29241\,
            I => \N__29238\
        );

    \I__5150\ : InMux
    port map (
            O => \N__29238\,
            I => \N__29235\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29235\,
            I => \N__29232\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__29232\,
            I => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\
        );

    \I__5147\ : CascadeMux
    port map (
            O => \N__29229\,
            I => \N__29226\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29226\,
            I => \N__29223\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__29223\,
            I => \N__29220\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__29220\,
            I => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\
        );

    \I__5143\ : InMux
    port map (
            O => \N__29217\,
            I => \N__29214\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__29214\,
            I => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29208\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29205\
        );

    \I__5139\ : Odrv4
    port map (
            O => \N__29205\,
            I => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29198\
        );

    \I__5137\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29195\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29198\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__29195\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__5134\ : CascadeMux
    port map (
            O => \N__29190\,
            I => \N__29187\
        );

    \I__5133\ : InMux
    port map (
            O => \N__29187\,
            I => \N__29184\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__29184\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29181\,
            I => \N__29178\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29178\,
            I => \N__29175\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__29175\,
            I => \N__29172\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__29172\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__29169\,
            I => \N__29166\
        );

    \I__5126\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29159\
        );

    \I__5124\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29156\
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__29159\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__29156\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__29148\,
            I => \N__29145\
        );

    \I__5119\ : Odrv12
    port map (
            O => \N__29145\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\
        );

    \I__5118\ : InMux
    port map (
            O => \N__29142\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_28\
        );

    \I__5117\ : InMux
    port map (
            O => \N__29139\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__5116\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29133\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29130\
        );

    \I__5114\ : Sp12to4
    port map (
            O => \N__29130\,
            I => \N__29127\
        );

    \I__5113\ : Span12Mux_v
    port map (
            O => \N__29127\,
            I => \N__29124\
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__29124\,
            I => \il_max_comp1_D1\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29118\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__29118\,
            I => \N__29115\
        );

    \I__5109\ : Odrv4
    port map (
            O => \N__29115\,
            I => \il_min_comp1_D1\
        );

    \I__5108\ : CascadeMux
    port map (
            O => \N__29112\,
            I => \N__29109\
        );

    \I__5107\ : InMux
    port map (
            O => \N__29109\,
            I => \N__29106\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__29106\,
            I => \N__29103\
        );

    \I__5105\ : Odrv12
    port map (
            O => \N__29103\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29097\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29097\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29091\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__29091\,
            I => \N__29088\
        );

    \I__5100\ : Sp12to4
    port map (
            O => \N__29088\,
            I => \N__29085\
        );

    \I__5099\ : Odrv12
    port map (
            O => \N__29085\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__29082\,
            I => \N__29079\
        );

    \I__5097\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29076\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29073\
        );

    \I__5095\ : Span4Mux_h
    port map (
            O => \N__29073\,
            I => \N__29070\
        );

    \I__5094\ : Odrv4
    port map (
            O => \N__29070\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__5093\ : InMux
    port map (
            O => \N__29067\,
            I => \N__29064\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__29064\,
            I => \N__29061\
        );

    \I__5091\ : Span4Mux_v
    port map (
            O => \N__29061\,
            I => \N__29058\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__29058\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__5089\ : CascadeMux
    port map (
            O => \N__29055\,
            I => \N__29052\
        );

    \I__5088\ : InMux
    port map (
            O => \N__29052\,
            I => \N__29049\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29046\
        );

    \I__5086\ : Span4Mux_v
    port map (
            O => \N__29046\,
            I => \N__29043\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__29043\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29040\,
            I => \N__29037\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__29037\,
            I => \N__29034\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__29034\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__29031\,
            I => \N__29028\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29028\,
            I => \N__29025\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__29025\,
            I => \N__29022\
        );

    \I__5078\ : Odrv12
    port map (
            O => \N__29022\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__5077\ : InMux
    port map (
            O => \N__29019\,
            I => \N__29016\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__29016\,
            I => \N__29013\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__29013\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__29010\,
            I => \N__29007\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29007\,
            I => \N__29004\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__29004\,
            I => \N__29001\
        );

    \I__5071\ : Span4Mux_h
    port map (
            O => \N__29001\,
            I => \N__28998\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__28998\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__5069\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28992\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__28992\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__5067\ : CascadeMux
    port map (
            O => \N__28989\,
            I => \N__28986\
        );

    \I__5066\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28983\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__28983\,
            I => \N__28980\
        );

    \I__5064\ : Odrv4
    port map (
            O => \N__28980\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__5063\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28974\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__28974\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__28971\,
            I => \N__28968\
        );

    \I__5060\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28965\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__28965\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__5058\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28959\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__28959\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__5056\ : CascadeMux
    port map (
            O => \N__28956\,
            I => \N__28953\
        );

    \I__5055\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28950\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__28950\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__5053\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28944\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28941\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__28941\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__5050\ : CascadeMux
    port map (
            O => \N__28938\,
            I => \N__28935\
        );

    \I__5049\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28932\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__28932\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__5047\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__5045\ : Span4Mux_v
    port map (
            O => \N__28923\,
            I => \N__28920\
        );

    \I__5044\ : Odrv4
    port map (
            O => \N__28920\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__5042\ : InMux
    port map (
            O => \N__28914\,
            I => \N__28911\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__28911\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__5040\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28905\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__28905\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__5038\ : CascadeMux
    port map (
            O => \N__28902\,
            I => \N__28899\
        );

    \I__5037\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28896\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__28896\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__5035\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28890\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__28890\,
            I => \N__28887\
        );

    \I__5033\ : Span4Mux_h
    port map (
            O => \N__28887\,
            I => \N__28884\
        );

    \I__5032\ : Odrv4
    port map (
            O => \N__28884\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__28881\,
            I => \N__28878\
        );

    \I__5030\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28875\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__28875\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__5028\ : InMux
    port map (
            O => \N__28872\,
            I => \N__28869\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__28869\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__28866\,
            I => \N__28863\
        );

    \I__5025\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28860\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__28860\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__5023\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28854\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__28854\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__28851\,
            I => \N__28848\
        );

    \I__5020\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28845\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__28845\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__5018\ : CascadeMux
    port map (
            O => \N__28842\,
            I => \N__28839\
        );

    \I__5017\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28836\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__28836\,
            I => \N__28833\
        );

    \I__5015\ : Odrv12
    port map (
            O => \N__28833\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__5014\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28827\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__28827\,
            I => \N__28824\
        );

    \I__5012\ : Odrv4
    port map (
            O => \N__28824\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__5011\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28818\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__28818\,
            I => \N__28815\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__28815\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__28812\,
            I => \N__28809\
        );

    \I__5007\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28806\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__28806\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__28803\,
            I => \N__28800\
        );

    \I__5004\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28794\
        );

    \I__5003\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28794\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__28794\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__5001\ : InMux
    port map (
            O => \N__28791\,
            I => \N__28788\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28785\
        );

    \I__4999\ : Span4Mux_h
    port map (
            O => \N__28785\,
            I => \N__28782\
        );

    \I__4998\ : Odrv4
    port map (
            O => \N__28782\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__28779\,
            I => \N__28776\
        );

    \I__4996\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28773\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__28773\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__4994\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28767\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__28767\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__4992\ : CascadeMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__4991\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__28758\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__4989\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28752\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__28752\,
            I => \N__28749\
        );

    \I__4987\ : Odrv12
    port map (
            O => \N__28749\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__4986\ : CascadeMux
    port map (
            O => \N__28746\,
            I => \N__28743\
        );

    \I__4985\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__28737\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__4982\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28731\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__28731\,
            I => \N__28728\
        );

    \I__4980\ : Odrv12
    port map (
            O => \N__28728\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__4979\ : CascadeMux
    port map (
            O => \N__28725\,
            I => \N__28722\
        );

    \I__4978\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__28719\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__4976\ : InMux
    port map (
            O => \N__28716\,
            I => \N__28713\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__28713\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__28710\,
            I => \N__28707\
        );

    \I__4973\ : InMux
    port map (
            O => \N__28707\,
            I => \N__28704\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__28704\,
            I => \N__28701\
        );

    \I__4971\ : Odrv4
    port map (
            O => \N__28701\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__4970\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28695\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__28695\,
            I => \N__28692\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__28689\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__28686\,
            I => \N__28683\
        );

    \I__4965\ : InMux
    port map (
            O => \N__28683\,
            I => \N__28680\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__28680\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__4963\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28671\
        );

    \I__4962\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28664\
        );

    \I__4961\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28664\
        );

    \I__4960\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28664\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__28671\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__28664\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__4957\ : InMux
    port map (
            O => \N__28659\,
            I => \N__28650\
        );

    \I__4956\ : InMux
    port map (
            O => \N__28658\,
            I => \N__28650\
        );

    \I__4955\ : InMux
    port map (
            O => \N__28657\,
            I => \N__28650\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__28650\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__28647\,
            I => \N__28642\
        );

    \I__4952\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28638\
        );

    \I__4951\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28631\
        );

    \I__4950\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28631\
        );

    \I__4949\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28631\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__28638\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__28631\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__28626\,
            I => \N__28622\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__28625\,
            I => \N__28618\
        );

    \I__4944\ : InMux
    port map (
            O => \N__28622\,
            I => \N__28611\
        );

    \I__4943\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28611\
        );

    \I__4942\ : InMux
    port map (
            O => \N__28618\,
            I => \N__28611\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__28611\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__4940\ : CascadeMux
    port map (
            O => \N__28608\,
            I => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\
        );

    \I__4939\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28596\
        );

    \I__4938\ : InMux
    port map (
            O => \N__28604\,
            I => \N__28596\
        );

    \I__4937\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28596\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__28596\,
            I => \N__28593\
        );

    \I__4935\ : Odrv4
    port map (
            O => \N__28593\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__4934\ : CascadeMux
    port map (
            O => \N__28590\,
            I => \N__28586\
        );

    \I__4933\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28578\
        );

    \I__4932\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28578\
        );

    \I__4931\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28578\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__28578\,
            I => \N__28575\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__28575\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__28572\,
            I => \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\
        );

    \I__4927\ : CascadeMux
    port map (
            O => \N__28569\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__4926\ : InMux
    port map (
            O => \N__28566\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__4925\ : CascadeMux
    port map (
            O => \N__28563\,
            I => \N__28559\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__28562\,
            I => \N__28556\
        );

    \I__4923\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28550\
        );

    \I__4922\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28550\
        );

    \I__4921\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28547\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__28550\,
            I => \N__28544\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__28547\,
            I => \N__28539\
        );

    \I__4918\ : Span4Mux_v
    port map (
            O => \N__28544\,
            I => \N__28539\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__28539\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__4916\ : InMux
    port map (
            O => \N__28536\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__4915\ : InMux
    port map (
            O => \N__28533\,
            I => \N__28528\
        );

    \I__4914\ : InMux
    port map (
            O => \N__28532\,
            I => \N__28523\
        );

    \I__4913\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28523\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__28528\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__28523\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__4910\ : InMux
    port map (
            O => \N__28518\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__4909\ : CascadeMux
    port map (
            O => \N__28515\,
            I => \N__28510\
        );

    \I__4908\ : InMux
    port map (
            O => \N__28514\,
            I => \N__28507\
        );

    \I__4907\ : InMux
    port map (
            O => \N__28513\,
            I => \N__28502\
        );

    \I__4906\ : InMux
    port map (
            O => \N__28510\,
            I => \N__28502\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__28507\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__28502\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__4903\ : InMux
    port map (
            O => \N__28497\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__4902\ : InMux
    port map (
            O => \N__28494\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__4901\ : InMux
    port map (
            O => \N__28491\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__4900\ : InMux
    port map (
            O => \N__28488\,
            I => \N__28483\
        );

    \I__4899\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28478\
        );

    \I__4898\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28478\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__28483\,
            I => \N__28474\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__28478\,
            I => \N__28471\
        );

    \I__4895\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28468\
        );

    \I__4894\ : Span4Mux_v
    port map (
            O => \N__28474\,
            I => \N__28461\
        );

    \I__4893\ : Span4Mux_v
    port map (
            O => \N__28471\,
            I => \N__28461\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__28468\,
            I => \N__28461\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__4890\ : Span4Mux_v
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__4889\ : Odrv4
    port map (
            O => \N__28455\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28452\,
            I => \N__28449\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__4886\ : Span4Mux_v
    port map (
            O => \N__28446\,
            I => \N__28441\
        );

    \I__4885\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28436\
        );

    \I__4884\ : InMux
    port map (
            O => \N__28444\,
            I => \N__28436\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__28441\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__28436\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__4881\ : InMux
    port map (
            O => \N__28431\,
            I => \N__28424\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28430\,
            I => \N__28424\
        );

    \I__4879\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28421\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28418\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28421\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__28418\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__4875\ : InMux
    port map (
            O => \N__28413\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__4874\ : CascadeMux
    port map (
            O => \N__28410\,
            I => \N__28407\
        );

    \I__4873\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28400\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28400\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28405\,
            I => \N__28397\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__28400\,
            I => \N__28394\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__28397\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4868\ : Odrv12
    port map (
            O => \N__28394\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4867\ : InMux
    port map (
            O => \N__28389\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__28386\,
            I => \N__28382\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__28385\,
            I => \N__28379\
        );

    \I__4864\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28376\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28373\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__28376\,
            I => \N__28367\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28367\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28364\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__28367\,
            I => \N__28361\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28364\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__28361\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__4856\ : InMux
    port map (
            O => \N__28356\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__4855\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28349\
        );

    \I__4854\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28345\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28349\,
            I => \N__28342\
        );

    \I__4852\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28339\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__28345\,
            I => \N__28336\
        );

    \I__4850\ : Span4Mux_h
    port map (
            O => \N__28342\,
            I => \N__28333\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__28339\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__28336\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4847\ : Odrv4
    port map (
            O => \N__28333\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__4846\ : InMux
    port map (
            O => \N__28326\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__28323\,
            I => \N__28319\
        );

    \I__4844\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28313\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28313\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28310\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28313\,
            I => \N__28307\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28310\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__28307\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28302\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__4837\ : CascadeMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__4836\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28291\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28288\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28285\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28291\,
            I => \N__28280\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28280\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__28285\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__28280\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__4829\ : InMux
    port map (
            O => \N__28275\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__4828\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28265\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28265\
        );

    \I__4826\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28262\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__28265\,
            I => \N__28259\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__28262\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4823\ : Odrv4
    port map (
            O => \N__28259\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28254\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__4821\ : CascadeMux
    port map (
            O => \N__28251\,
            I => \N__28247\
        );

    \I__4820\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28241\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28247\,
            I => \N__28241\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28246\,
            I => \N__28238\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28241\,
            I => \N__28235\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__28238\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4815\ : Odrv4
    port map (
            O => \N__28235\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28230\,
            I => \bfn_11_8_0_\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28227\,
            I => \N__28220\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28226\,
            I => \N__28220\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28225\,
            I => \N__28217\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28214\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28217\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4808\ : Odrv4
    port map (
            O => \N__28214\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28209\,
            I => \bfn_11_6_0_\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28206\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28203\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__4804\ : InMux
    port map (
            O => \N__28200\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__4803\ : InMux
    port map (
            O => \N__28197\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28194\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28191\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28181\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28187\,
            I => \N__28181\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28186\,
            I => \N__28178\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__28181\,
            I => \N__28175\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__28178\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__28175\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28170\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__28167\,
            I => \N__28162\
        );

    \I__4792\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28159\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28154\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28154\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__28159\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28154\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__4787\ : InMux
    port map (
            O => \N__28149\,
            I => \bfn_11_7_0_\
        );

    \I__4786\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \N__28143\
        );

    \I__4785\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28136\
        );

    \I__4784\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28136\
        );

    \I__4783\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28133\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__28136\,
            I => \N__28130\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__28133\,
            I => \N__28125\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__28130\,
            I => \N__28125\
        );

    \I__4779\ : Span4Mux_v
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__4778\ : Span4Mux_v
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__4777\ : Odrv4
    port map (
            O => \N__28119\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__4776\ : InMux
    port map (
            O => \N__28116\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__4775\ : InMux
    port map (
            O => \N__28113\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__4774\ : InMux
    port map (
            O => \N__28110\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__4773\ : InMux
    port map (
            O => \N__28107\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28104\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__4771\ : InMux
    port map (
            O => \N__28101\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28098\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__4769\ : CascadeMux
    port map (
            O => \N__28095\,
            I => \N__28092\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28089\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__28086\,
            I => \N__28083\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__4764\ : Span4Mux_h
    port map (
            O => \N__28080\,
            I => \N__28077\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__28077\,
            I => \N__28074\
        );

    \I__4762\ : Odrv4
    port map (
            O => \N__28074\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28068\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__28068\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28065\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__4758\ : CascadeMux
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28056\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__28056\,
            I => \N__28053\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__28053\,
            I => \N__28050\
        );

    \I__4754\ : Sp12to4
    port map (
            O => \N__28050\,
            I => \N__28047\
        );

    \I__4753\ : Span12Mux_h
    port map (
            O => \N__28047\,
            I => \N__28044\
        );

    \I__4752\ : Odrv12
    port map (
            O => \N__28044\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__4751\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28038\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__28038\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28035\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__28032\,
            I => \N__28029\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28029\,
            I => \N__28026\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__28026\,
            I => \N__28023\
        );

    \I__4745\ : Span12Mux_h
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__4744\ : Span12Mux_h
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__4743\ : Odrv12
    port map (
            O => \N__28017\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__4742\ : InMux
    port map (
            O => \N__28014\,
            I => \N__28011\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__28011\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__4740\ : InMux
    port map (
            O => \N__28008\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27999\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__27999\,
            I => \N__27996\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__27996\,
            I => \N__27993\
        );

    \I__4735\ : Sp12to4
    port map (
            O => \N__27993\,
            I => \N__27990\
        );

    \I__4734\ : Span12Mux_h
    port map (
            O => \N__27990\,
            I => \N__27987\
        );

    \I__4733\ : Odrv12
    port map (
            O => \N__27987\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__4732\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__27981\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__4730\ : InMux
    port map (
            O => \N__27978\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__4729\ : CascadeMux
    port map (
            O => \N__27975\,
            I => \N__27972\
        );

    \I__4728\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27969\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27966\
        );

    \I__4726\ : Span4Mux_v
    port map (
            O => \N__27966\,
            I => \N__27963\
        );

    \I__4725\ : Sp12to4
    port map (
            O => \N__27963\,
            I => \N__27960\
        );

    \I__4724\ : Span12Mux_h
    port map (
            O => \N__27960\,
            I => \N__27957\
        );

    \I__4723\ : Odrv12
    port map (
            O => \N__27957\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__4722\ : InMux
    port map (
            O => \N__27954\,
            I => \N__27951\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__27951\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__4720\ : InMux
    port map (
            O => \N__27948\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__4719\ : CascadeMux
    port map (
            O => \N__27945\,
            I => \N__27942\
        );

    \I__4718\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27939\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27936\
        );

    \I__4716\ : Span4Mux_v
    port map (
            O => \N__27936\,
            I => \N__27933\
        );

    \I__4715\ : Span4Mux_h
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__4714\ : Sp12to4
    port map (
            O => \N__27930\,
            I => \N__27927\
        );

    \I__4713\ : Odrv12
    port map (
            O => \N__27927\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__4712\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27921\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__27921\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__4710\ : InMux
    port map (
            O => \N__27918\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__4709\ : InMux
    port map (
            O => \N__27915\,
            I => \N__27903\
        );

    \I__4708\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27903\
        );

    \I__4707\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27896\
        );

    \I__4706\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27896\
        );

    \I__4705\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27896\
        );

    \I__4704\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27889\
        );

    \I__4703\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27889\
        );

    \I__4702\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27889\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__27903\,
            I => \N__27886\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27881\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__27889\,
            I => \N__27881\
        );

    \I__4698\ : Span12Mux_h
    port map (
            O => \N__27886\,
            I => \N__27878\
        );

    \I__4697\ : Span12Mux_h
    port map (
            O => \N__27881\,
            I => \N__27875\
        );

    \I__4696\ : Odrv12
    port map (
            O => \N__27878\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__4695\ : Odrv12
    port map (
            O => \N__27875\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__27870\,
            I => \N__27867\
        );

    \I__4693\ : InMux
    port map (
            O => \N__27867\,
            I => \N__27864\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__27864\,
            I => \N__27861\
        );

    \I__4691\ : Odrv12
    port map (
            O => \N__27861\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__4690\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27855\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__27855\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__4688\ : InMux
    port map (
            O => \N__27852\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__4687\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__27846\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__4685\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27840\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__27840\,
            I => \N__27837\
        );

    \I__4683\ : Odrv12
    port map (
            O => \N__27837\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__4682\ : InMux
    port map (
            O => \N__27834\,
            I => \bfn_10_28_0_\
        );

    \I__4681\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27828\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27825\
        );

    \I__4679\ : Span4Mux_v
    port map (
            O => \N__27825\,
            I => \N__27822\
        );

    \I__4678\ : Sp12to4
    port map (
            O => \N__27822\,
            I => \N__27819\
        );

    \I__4677\ : Span12Mux_h
    port map (
            O => \N__27819\,
            I => \N__27816\
        );

    \I__4676\ : Odrv12
    port map (
            O => \N__27816\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__4674\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27807\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__27807\,
            I => \N__27804\
        );

    \I__4672\ : Span12Mux_h
    port map (
            O => \N__27804\,
            I => \N__27801\
        );

    \I__4671\ : Odrv12
    port map (
            O => \N__27801\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__4670\ : InMux
    port map (
            O => \N__27798\,
            I => \N__27795\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__27795\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__4668\ : InMux
    port map (
            O => \N__27792\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__4667\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27786\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__27786\,
            I => \N__27783\
        );

    \I__4665\ : Span12Mux_h
    port map (
            O => \N__27783\,
            I => \N__27780\
        );

    \I__4664\ : Span12Mux_h
    port map (
            O => \N__27780\,
            I => \N__27777\
        );

    \I__4663\ : Odrv12
    port map (
            O => \N__27777\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__4662\ : CascadeMux
    port map (
            O => \N__27774\,
            I => \N__27771\
        );

    \I__4661\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27768\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__4659\ : Span4Mux_h
    port map (
            O => \N__27765\,
            I => \N__27762\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__27762\,
            I => \N__27759\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__27759\,
            I => \N__27756\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__27756\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__27753\,
            I => \N__27750\
        );

    \I__4654\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27747\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__27747\,
            I => \N__27744\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__27744\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__4651\ : InMux
    port map (
            O => \N__27741\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__4650\ : InMux
    port map (
            O => \N__27738\,
            I => \N__27735\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27732\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__27732\,
            I => \N__27729\
        );

    \I__4647\ : Sp12to4
    port map (
            O => \N__27729\,
            I => \N__27726\
        );

    \I__4646\ : Span12Mux_h
    port map (
            O => \N__27726\,
            I => \N__27723\
        );

    \I__4645\ : Odrv12
    port map (
            O => \N__27723\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__27720\,
            I => \N__27717\
        );

    \I__4643\ : InMux
    port map (
            O => \N__27717\,
            I => \N__27714\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__27714\,
            I => \N__27711\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__27711\,
            I => \N__27708\
        );

    \I__4640\ : Span4Mux_h
    port map (
            O => \N__27708\,
            I => \N__27705\
        );

    \I__4639\ : Span4Mux_h
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__27702\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__4637\ : InMux
    port map (
            O => \N__27699\,
            I => \N__27696\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__27696\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__4635\ : InMux
    port map (
            O => \N__27693\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__4634\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27687\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__4631\ : Sp12to4
    port map (
            O => \N__27681\,
            I => \N__27678\
        );

    \I__4630\ : Span12Mux_h
    port map (
            O => \N__27678\,
            I => \N__27675\
        );

    \I__4629\ : Odrv12
    port map (
            O => \N__27675\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__4627\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27666\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__27666\,
            I => \N__27663\
        );

    \I__4625\ : Span4Mux_v
    port map (
            O => \N__27663\,
            I => \N__27660\
        );

    \I__4624\ : Span4Mux_h
    port map (
            O => \N__27660\,
            I => \N__27657\
        );

    \I__4623\ : Span4Mux_h
    port map (
            O => \N__27657\,
            I => \N__27654\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__27654\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__4621\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27648\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__27648\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__4619\ : InMux
    port map (
            O => \N__27645\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__4618\ : InMux
    port map (
            O => \N__27642\,
            I => \N__27639\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__27639\,
            I => \N__27636\
        );

    \I__4616\ : Span4Mux_v
    port map (
            O => \N__27636\,
            I => \N__27633\
        );

    \I__4615\ : Span4Mux_h
    port map (
            O => \N__27633\,
            I => \N__27630\
        );

    \I__4614\ : Sp12to4
    port map (
            O => \N__27630\,
            I => \N__27627\
        );

    \I__4613\ : Odrv12
    port map (
            O => \N__27627\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__27624\,
            I => \N__27621\
        );

    \I__4611\ : InMux
    port map (
            O => \N__27621\,
            I => \N__27618\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__27618\,
            I => \N__27615\
        );

    \I__4609\ : Sp12to4
    port map (
            O => \N__27615\,
            I => \N__27612\
        );

    \I__4608\ : Span12Mux_s5_v
    port map (
            O => \N__27612\,
            I => \N__27609\
        );

    \I__4607\ : Odrv12
    port map (
            O => \N__27609\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__4606\ : InMux
    port map (
            O => \N__27606\,
            I => \N__27603\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__27603\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__4604\ : InMux
    port map (
            O => \N__27600\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__4603\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27594\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__27594\,
            I => \N__27591\
        );

    \I__4601\ : Span12Mux_s5_v
    port map (
            O => \N__27591\,
            I => \N__27588\
        );

    \I__4600\ : Odrv12
    port map (
            O => \N__27588\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__27585\,
            I => \N__27582\
        );

    \I__4598\ : InMux
    port map (
            O => \N__27582\,
            I => \N__27579\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__27579\,
            I => \N__27576\
        );

    \I__4596\ : Span12Mux_s7_v
    port map (
            O => \N__27576\,
            I => \N__27573\
        );

    \I__4595\ : Span12Mux_h
    port map (
            O => \N__27573\,
            I => \N__27570\
        );

    \I__4594\ : Odrv12
    port map (
            O => \N__27570\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__4593\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27564\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__27564\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__4591\ : InMux
    port map (
            O => \N__27561\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__4590\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27555\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__27555\,
            I => \N__27552\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__27552\,
            I => \N__27549\
        );

    \I__4587\ : Sp12to4
    port map (
            O => \N__27549\,
            I => \N__27546\
        );

    \I__4586\ : Odrv12
    port map (
            O => \N__27546\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__27543\,
            I => \N__27540\
        );

    \I__4584\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27537\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__27537\,
            I => \N__27534\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__27534\,
            I => \N__27531\
        );

    \I__4581\ : Sp12to4
    port map (
            O => \N__27531\,
            I => \N__27528\
        );

    \I__4580\ : Span12Mux_h
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__4579\ : Odrv12
    port map (
            O => \N__27525\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__4578\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27519\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__27519\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__4576\ : InMux
    port map (
            O => \N__27516\,
            I => \bfn_10_27_0_\
        );

    \I__4575\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27510\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__27510\,
            I => \N__27507\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__27501\,
            I => \N__27498\
        );

    \I__4570\ : Odrv4
    port map (
            O => \N__27498\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__4569\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27489\
        );

    \I__4568\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27489\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__4566\ : Span12Mux_v
    port map (
            O => \N__27486\,
            I => \N__27483\
        );

    \I__4565\ : Span12Mux_h
    port map (
            O => \N__27483\,
            I => \N__27480\
        );

    \I__4564\ : Odrv12
    port map (
            O => \N__27480\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27474\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__27474\,
            I => \N__27471\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__4560\ : Sp12to4
    port map (
            O => \N__27468\,
            I => \N__27465\
        );

    \I__4559\ : Span12Mux_h
    port map (
            O => \N__27465\,
            I => \N__27462\
        );

    \I__4558\ : Odrv12
    port map (
            O => \N__27462\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__4557\ : InMux
    port map (
            O => \N__27459\,
            I => \N__27456\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__27453\,
            I => \N__27450\
        );

    \I__4554\ : Odrv4
    port map (
            O => \N__27450\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__4553\ : InMux
    port map (
            O => \N__27447\,
            I => \N__27443\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27446\,
            I => \N__27440\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__27443\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__27440\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__27432\,
            I => \N__27428\
        );

    \I__4547\ : InMux
    port map (
            O => \N__27431\,
            I => \N__27424\
        );

    \I__4546\ : Span4Mux_h
    port map (
            O => \N__27428\,
            I => \N__27421\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27427\,
            I => \N__27418\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__27424\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__27421\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__27418\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27408\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__4539\ : Span4Mux_h
    port map (
            O => \N__27405\,
            I => \N__27402\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__27402\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__27399\,
            I => \N__27396\
        );

    \I__4536\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27393\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__27393\,
            I => \N__27389\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27385\
        );

    \I__4533\ : Span4Mux_v
    port map (
            O => \N__27389\,
            I => \N__27382\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27379\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__27385\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__27382\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__27379\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27372\,
            I => \N__27368\
        );

    \I__4527\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27365\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27368\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27365\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__4524\ : InMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__27357\,
            I => \N__27354\
        );

    \I__4522\ : Span4Mux_h
    port map (
            O => \N__27354\,
            I => \N__27351\
        );

    \I__4521\ : Odrv4
    port map (
            O => \N__27351\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4519\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27341\
        );

    \I__4518\ : InMux
    port map (
            O => \N__27344\,
            I => \N__27338\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27341\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__27338\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27326\
        );

    \I__4513\ : InMux
    port map (
            O => \N__27329\,
            I => \N__27322\
        );

    \I__4512\ : Span4Mux_h
    port map (
            O => \N__27326\,
            I => \N__27319\
        );

    \I__4511\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27316\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__27322\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__27319\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__27316\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27304\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27308\,
            I => \N__27301\
        );

    \I__4505\ : InMux
    port map (
            O => \N__27307\,
            I => \N__27298\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__27304\,
            I => \N__27295\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__27301\,
            I => \N__27292\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__27298\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__4501\ : Odrv12
    port map (
            O => \N__27295\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__27292\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__4499\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__27279\,
            I => \N__27276\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__27276\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27270\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27266\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27263\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__27266\,
            I => \N__27258\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__27263\,
            I => \N__27258\
        );

    \I__4490\ : Span4Mux_h
    port map (
            O => \N__27258\,
            I => \N__27255\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__4488\ : Odrv4
    port map (
            O => \N__27252\,
            I => \pwm_generator_inst.O_10\
        );

    \I__4487\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27245\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27242\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__27245\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__27242\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4482\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27231\,
            I => \N__27227\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27223\
        );

    \I__4479\ : Span4Mux_h
    port map (
            O => \N__27227\,
            I => \N__27220\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27217\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__27223\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__4476\ : Odrv4
    port map (
            O => \N__27220\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27217\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__4474\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__27207\,
            I => \N__27204\
        );

    \I__4472\ : Span4Mux_h
    port map (
            O => \N__27204\,
            I => \N__27201\
        );

    \I__4471\ : Odrv4
    port map (
            O => \N__27201\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27198\,
            I => \N__27195\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__4468\ : Span4Mux_v
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__4467\ : Sp12to4
    port map (
            O => \N__27189\,
            I => \N__27186\
        );

    \I__4466\ : Span12Mux_h
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4465\ : Odrv12
    port map (
            O => \N__27183\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__27180\,
            I => \N__27177\
        );

    \I__4463\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__27171\,
            I => \N__27168\
        );

    \I__4460\ : Span4Mux_h
    port map (
            O => \N__27168\,
            I => \N__27165\
        );

    \I__4459\ : Span4Mux_h
    port map (
            O => \N__27165\,
            I => \N__27162\
        );

    \I__4458\ : Odrv4
    port map (
            O => \N__27162\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27156\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__4455\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__27150\,
            I => \N__27147\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__4452\ : Sp12to4
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__4451\ : Span12Mux_h
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__4450\ : Odrv12
    port map (
            O => \N__27138\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27129\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__27126\,
            I => \N__27123\
        );

    \I__4445\ : Span4Mux_h
    port map (
            O => \N__27123\,
            I => \N__27120\
        );

    \I__4444\ : Span4Mux_h
    port map (
            O => \N__27120\,
            I => \N__27117\
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__27117\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__27114\,
            I => \N__27111\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27111\,
            I => \N__27108\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__27108\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__4439\ : InMux
    port map (
            O => \N__27105\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27098\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27094\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27091\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27088\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27094\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4433\ : Odrv12
    port map (
            O => \N__27091\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__27088\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27075\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__27080\,
            I => \N__27072\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27079\,
            I => \N__27069\
        );

    \I__4428\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27066\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__27075\,
            I => \N__27063\
        );

    \I__4426\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27060\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__27069\,
            I => \N__27057\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__27066\,
            I => \N__27054\
        );

    \I__4423\ : Span4Mux_h
    port map (
            O => \N__27063\,
            I => \N__27051\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27060\,
            I => \N__27048\
        );

    \I__4421\ : Span12Mux_s11_v
    port map (
            O => \N__27057\,
            I => \N__27045\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__27054\,
            I => \N__27038\
        );

    \I__4419\ : Span4Mux_v
    port map (
            O => \N__27051\,
            I => \N__27038\
        );

    \I__4418\ : Span4Mux_h
    port map (
            O => \N__27048\,
            I => \N__27038\
        );

    \I__4417\ : Odrv12
    port map (
            O => \N__27045\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__27038\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__27033\,
            I => \N__27030\
        );

    \I__4414\ : InMux
    port map (
            O => \N__27030\,
            I => \N__27024\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27029\,
            I => \N__27024\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__27024\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__4411\ : CEMux
    port map (
            O => \N__27021\,
            I => \N__27000\
        );

    \I__4410\ : CEMux
    port map (
            O => \N__27020\,
            I => \N__27000\
        );

    \I__4409\ : CEMux
    port map (
            O => \N__27019\,
            I => \N__27000\
        );

    \I__4408\ : CEMux
    port map (
            O => \N__27018\,
            I => \N__27000\
        );

    \I__4407\ : CEMux
    port map (
            O => \N__27017\,
            I => \N__27000\
        );

    \I__4406\ : CEMux
    port map (
            O => \N__27016\,
            I => \N__27000\
        );

    \I__4405\ : CEMux
    port map (
            O => \N__27015\,
            I => \N__27000\
        );

    \I__4404\ : GlobalMux
    port map (
            O => \N__27000\,
            I => \N__26997\
        );

    \I__4403\ : gio2CtrlBuf
    port map (
            O => \N__26997\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__4402\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26990\
        );

    \I__4401\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26987\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26984\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__26987\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__26984\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__4397\ : InMux
    port map (
            O => \N__26979\,
            I => \N__26975\
        );

    \I__4396\ : InMux
    port map (
            O => \N__26978\,
            I => \N__26972\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__26975\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__26972\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__4393\ : InMux
    port map (
            O => \N__26967\,
            I => \N__26961\
        );

    \I__4392\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26954\
        );

    \I__4391\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26954\
        );

    \I__4390\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26954\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__26961\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__26954\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__4387\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26946\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__26946\,
            I => \N__26943\
        );

    \I__4385\ : Span4Mux_h
    port map (
            O => \N__26943\,
            I => \N__26940\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__26940\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__4383\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__4381\ : Span4Mux_h
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__26928\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__4379\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__26922\,
            I => \N__26919\
        );

    \I__4377\ : Span4Mux_h
    port map (
            O => \N__26919\,
            I => \N__26916\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__26916\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__4375\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26905\
        );

    \I__4374\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26893\
        );

    \I__4373\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26893\
        );

    \I__4372\ : InMux
    port map (
            O => \N__26910\,
            I => \N__26893\
        );

    \I__4371\ : InMux
    port map (
            O => \N__26909\,
            I => \N__26893\
        );

    \I__4370\ : InMux
    port map (
            O => \N__26908\,
            I => \N__26890\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__26905\,
            I => \N__26887\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__26904\,
            I => \N__26883\
        );

    \I__4367\ : InMux
    port map (
            O => \N__26903\,
            I => \N__26878\
        );

    \I__4366\ : InMux
    port map (
            O => \N__26902\,
            I => \N__26878\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__26893\,
            I => \N__26873\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__26890\,
            I => \N__26873\
        );

    \I__4363\ : Span4Mux_h
    port map (
            O => \N__26887\,
            I => \N__26870\
        );

    \I__4362\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26865\
        );

    \I__4361\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26865\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__26878\,
            I => \N__26862\
        );

    \I__4359\ : Span4Mux_v
    port map (
            O => \N__26873\,
            I => \N__26859\
        );

    \I__4358\ : Span4Mux_h
    port map (
            O => \N__26870\,
            I => \N__26854\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__26865\,
            I => \N__26854\
        );

    \I__4356\ : Span4Mux_h
    port map (
            O => \N__26862\,
            I => \N__26851\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__26859\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__26854\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__4353\ : Odrv4
    port map (
            O => \N__26851\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__4352\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26838\
        );

    \I__4351\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26838\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__26838\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__4349\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26832\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__26832\,
            I => \N__26828\
        );

    \I__4347\ : InMux
    port map (
            O => \N__26831\,
            I => \N__26824\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__26828\,
            I => \N__26821\
        );

    \I__4345\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26818\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__26824\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__26821\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__26818\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__4341\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26808\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__26808\,
            I => \N__26802\
        );

    \I__4339\ : InMux
    port map (
            O => \N__26807\,
            I => \N__26799\
        );

    \I__4338\ : InMux
    port map (
            O => \N__26806\,
            I => \N__26794\
        );

    \I__4337\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26794\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__26802\,
            I => \N__26789\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26789\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__26794\,
            I => \N__26786\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__26789\,
            I => \N__26783\
        );

    \I__4332\ : Span4Mux_h
    port map (
            O => \N__26786\,
            I => \N__26780\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__26783\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__4330\ : Odrv4
    port map (
            O => \N__26780\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__26775\,
            I => \N__26772\
        );

    \I__4328\ : InMux
    port map (
            O => \N__26772\,
            I => \N__26766\
        );

    \I__4327\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26766\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__26766\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__4325\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26759\
        );

    \I__4324\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26755\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__26759\,
            I => \N__26752\
        );

    \I__4322\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26749\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__26755\,
            I => \N__26745\
        );

    \I__4320\ : Span4Mux_h
    port map (
            O => \N__26752\,
            I => \N__26742\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26739\
        );

    \I__4318\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26736\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__26745\,
            I => \N__26733\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__26742\,
            I => \N__26730\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__26739\,
            I => \N__26725\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26725\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__26733\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__26730\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__4311\ : Odrv4
    port map (
            O => \N__26725\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__4310\ : InMux
    port map (
            O => \N__26718\,
            I => \N__26713\
        );

    \I__4309\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26710\
        );

    \I__4308\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26707\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__26713\,
            I => \N__26704\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__26710\,
            I => \N__26701\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__26707\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__4304\ : Odrv12
    port map (
            O => \N__26704\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__26701\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__4302\ : InMux
    port map (
            O => \N__26694\,
            I => \N__26688\
        );

    \I__4301\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26688\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__26688\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__26685\,
            I => \N__26682\
        );

    \I__4298\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26679\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__26679\,
            I => \N__26675\
        );

    \I__4296\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26672\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__26675\,
            I => \N__26669\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__26672\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__26669\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__26664\,
            I => \N__26658\
        );

    \I__4291\ : InMux
    port map (
            O => \N__26663\,
            I => \N__26653\
        );

    \I__4290\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26653\
        );

    \I__4289\ : InMux
    port map (
            O => \N__26661\,
            I => \N__26650\
        );

    \I__4288\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26647\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__26653\,
            I => \N__26644\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__26650\,
            I => \N__26639\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__26647\,
            I => \N__26639\
        );

    \I__4284\ : Span4Mux_h
    port map (
            O => \N__26644\,
            I => \N__26636\
        );

    \I__4283\ : Span4Mux_v
    port map (
            O => \N__26639\,
            I => \N__26633\
        );

    \I__4282\ : Odrv4
    port map (
            O => \N__26636\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__26633\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__26628\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\
        );

    \I__4279\ : InMux
    port map (
            O => \N__26625\,
            I => \N__26620\
        );

    \I__4278\ : InMux
    port map (
            O => \N__26624\,
            I => \N__26617\
        );

    \I__4277\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26614\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__26620\,
            I => \N__26611\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__26617\,
            I => \N__26608\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__26614\,
            I => \N__26603\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__26611\,
            I => \N__26603\
        );

    \I__4272\ : Span4Mux_v
    port map (
            O => \N__26608\,
            I => \N__26600\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__26603\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__26600\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__4269\ : InMux
    port map (
            O => \N__26595\,
            I => \N__26591\
        );

    \I__4268\ : InMux
    port map (
            O => \N__26594\,
            I => \N__26587\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26584\
        );

    \I__4266\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26581\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__26587\,
            I => \N__26575\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__26584\,
            I => \N__26575\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__26581\,
            I => \N__26572\
        );

    \I__4262\ : InMux
    port map (
            O => \N__26580\,
            I => \N__26569\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__26575\,
            I => \N__26566\
        );

    \I__4260\ : Span4Mux_v
    port map (
            O => \N__26572\,
            I => \N__26561\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__26569\,
            I => \N__26561\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__26566\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__26561\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__4256\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26550\
        );

    \I__4255\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26550\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__26550\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__4253\ : InMux
    port map (
            O => \N__26547\,
            I => \N__26544\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__26544\,
            I => \N__26540\
        );

    \I__4251\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26536\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__26540\,
            I => \N__26533\
        );

    \I__4249\ : InMux
    port map (
            O => \N__26539\,
            I => \N__26530\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__26536\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__26533\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__26530\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__4245\ : CascadeMux
    port map (
            O => \N__26523\,
            I => \N__26518\
        );

    \I__4244\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26515\
        );

    \I__4243\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26511\
        );

    \I__4242\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26508\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__26515\,
            I => \N__26505\
        );

    \I__4240\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26502\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__26511\,
            I => \N__26499\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__26508\,
            I => \N__26496\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__26505\,
            I => \N__26493\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26490\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__26499\,
            I => \N__26487\
        );

    \I__4234\ : Span4Mux_v
    port map (
            O => \N__26496\,
            I => \N__26484\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__26493\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__26490\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__26487\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__26484\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__26475\,
            I => \N__26472\
        );

    \I__4228\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26466\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26471\,
            I => \N__26466\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__26466\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__4225\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26460\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__26460\,
            I => \N__26455\
        );

    \I__4223\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26452\
        );

    \I__4222\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26449\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__26455\,
            I => \N__26446\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26443\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__26449\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__4218\ : Odrv4
    port map (
            O => \N__26446\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__4217\ : Odrv12
    port map (
            O => \N__26443\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__4216\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26432\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26429\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__26432\,
            I => \N__26426\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__26429\,
            I => \N__26419\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__26426\,
            I => \N__26419\
        );

    \I__4211\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26414\
        );

    \I__4210\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26414\
        );

    \I__4209\ : Span4Mux_v
    port map (
            O => \N__26419\,
            I => \N__26409\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__26414\,
            I => \N__26409\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__26409\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26402\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26399\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__26402\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__26399\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__26394\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26383\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26390\,
            I => \N__26383\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26378\
        );

    \I__4198\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26378\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26383\,
            I => \N__26375\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26378\,
            I => \N__26372\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__26375\,
            I => \N__26369\
        );

    \I__4194\ : Odrv4
    port map (
            O => \N__26372\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__4193\ : Odrv4
    port map (
            O => \N__26369\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26360\
        );

    \I__4191\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26357\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26360\,
            I => \N__26352\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26357\,
            I => \N__26349\
        );

    \I__4188\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26346\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26343\
        );

    \I__4186\ : Span4Mux_h
    port map (
            O => \N__26352\,
            I => \N__26340\
        );

    \I__4185\ : Span4Mux_v
    port map (
            O => \N__26349\,
            I => \N__26335\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__26346\,
            I => \N__26335\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__26343\,
            I => \N__26332\
        );

    \I__4182\ : Span4Mux_v
    port map (
            O => \N__26340\,
            I => \N__26327\
        );

    \I__4181\ : Span4Mux_h
    port map (
            O => \N__26335\,
            I => \N__26327\
        );

    \I__4180\ : Span4Mux_v
    port map (
            O => \N__26332\,
            I => \N__26324\
        );

    \I__4179\ : Odrv4
    port map (
            O => \N__26327\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4178\ : Odrv4
    port map (
            O => \N__26324\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__4177\ : InMux
    port map (
            O => \N__26319\,
            I => \N__26316\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__26316\,
            I => \N__26313\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__26313\,
            I => \N__26308\
        );

    \I__4174\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26305\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26302\
        );

    \I__4172\ : Span4Mux_v
    port map (
            O => \N__26308\,
            I => \N__26299\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__26305\,
            I => \N__26296\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__26302\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__26299\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__26296\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26283\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26278\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26287\,
            I => \N__26278\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26275\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__26283\,
            I => \N__26272\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__26278\,
            I => \N__26269\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__26275\,
            I => \N__26266\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__26272\,
            I => \N__26261\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__26269\,
            I => \N__26261\
        );

    \I__4158\ : Span4Mux_h
    port map (
            O => \N__26266\,
            I => \N__26258\
        );

    \I__4157\ : Odrv4
    port map (
            O => \N__26261\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__26258\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26247\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26252\,
            I => \N__26247\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__26247\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26244\,
            I => \N__26240\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26236\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__26240\,
            I => \N__26233\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26230\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26236\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4147\ : Odrv12
    port map (
            O => \N__26233\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__26230\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__4145\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26219\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26214\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__26219\,
            I => \N__26211\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26218\,
            I => \N__26208\
        );

    \I__4141\ : InMux
    port map (
            O => \N__26217\,
            I => \N__26205\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__26214\,
            I => \N__26202\
        );

    \I__4139\ : Span4Mux_v
    port map (
            O => \N__26211\,
            I => \N__26195\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__26208\,
            I => \N__26195\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__26205\,
            I => \N__26195\
        );

    \I__4136\ : Span4Mux_h
    port map (
            O => \N__26202\,
            I => \N__26190\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__26195\,
            I => \N__26190\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__26190\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26181\
        );

    \I__4132\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26181\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__26181\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__4130\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26171\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26177\,
            I => \N__26171\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26167\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26164\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26170\,
            I => \N__26161\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__26167\,
            I => \N__26156\
        );

    \I__4124\ : Span4Mux_v
    port map (
            O => \N__26164\,
            I => \N__26156\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26153\
        );

    \I__4122\ : Span4Mux_v
    port map (
            O => \N__26156\,
            I => \N__26150\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__26153\,
            I => \N__26147\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__26150\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__26147\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__4118\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26139\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__26139\,
            I => \N__26135\
        );

    \I__4116\ : InMux
    port map (
            O => \N__26138\,
            I => \N__26132\
        );

    \I__4115\ : Odrv4
    port map (
            O => \N__26135\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__26132\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__26127\,
            I => \N__26124\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26118\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26118\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__26118\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__4109\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26111\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26108\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26105\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__26108\,
            I => \N__26098\
        );

    \I__4105\ : Span4Mux_v
    port map (
            O => \N__26105\,
            I => \N__26098\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26104\,
            I => \N__26095\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26103\,
            I => \N__26092\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__26098\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26095\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26092\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__4099\ : InMux
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__26082\,
            I => \N__26077\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26081\,
            I => \N__26074\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26080\,
            I => \N__26071\
        );

    \I__4095\ : Span4Mux_h
    port map (
            O => \N__26077\,
            I => \N__26068\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26074\,
            I => \N__26065\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__26071\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__26068\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4091\ : Odrv12
    port map (
            O => \N__26065\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26058\,
            I => \N__26053\
        );

    \I__4089\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26050\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26056\,
            I => \N__26047\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26053\,
            I => \N__26043\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__26040\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__26047\,
            I => \N__26037\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26046\,
            I => \N__26034\
        );

    \I__4083\ : Span4Mux_v
    port map (
            O => \N__26043\,
            I => \N__26031\
        );

    \I__4082\ : Span4Mux_v
    port map (
            O => \N__26040\,
            I => \N__26028\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__26037\,
            I => \N__26025\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__26034\,
            I => \N__26022\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__26031\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__26028\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__26025\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__26022\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26009\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26005\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26009\,
            I => \N__26002\
        );

    \I__4072\ : InMux
    port map (
            O => \N__26008\,
            I => \N__25999\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__26005\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__26002\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__25999\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__4068\ : InMux
    port map (
            O => \N__25992\,
            I => \N__25989\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__25989\,
            I => \N__25986\
        );

    \I__4066\ : Odrv12
    port map (
            O => \N__25986\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__4065\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25978\
        );

    \I__4064\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25974\
        );

    \I__4063\ : InMux
    port map (
            O => \N__25981\,
            I => \N__25971\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__25978\,
            I => \N__25968\
        );

    \I__4061\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25965\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__25974\,
            I => \N__25962\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__25971\,
            I => \N__25957\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__25968\,
            I => \N__25957\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25954\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__25962\,
            I => \N__25947\
        );

    \I__4055\ : Span4Mux_v
    port map (
            O => \N__25957\,
            I => \N__25947\
        );

    \I__4054\ : Span4Mux_v
    port map (
            O => \N__25954\,
            I => \N__25947\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__25947\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__4052\ : InMux
    port map (
            O => \N__25944\,
            I => \N__25941\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__25941\,
            I => \N__25938\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__25938\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\
        );

    \I__4049\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25932\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__25932\,
            I => \N__25929\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__25929\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__25926\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23_cascade_\
        );

    \I__4045\ : InMux
    port map (
            O => \N__25923\,
            I => \N__25920\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__25920\,
            I => \N__25917\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__25917\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__25914\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__4041\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25908\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__25908\,
            I => \N__25903\
        );

    \I__4039\ : InMux
    port map (
            O => \N__25907\,
            I => \N__25900\
        );

    \I__4038\ : InMux
    port map (
            O => \N__25906\,
            I => \N__25897\
        );

    \I__4037\ : Span4Mux_v
    port map (
            O => \N__25903\,
            I => \N__25894\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25891\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__25897\,
            I => \N__25886\
        );

    \I__4034\ : Span4Mux_v
    port map (
            O => \N__25894\,
            I => \N__25886\
        );

    \I__4033\ : Span4Mux_h
    port map (
            O => \N__25891\,
            I => \N__25883\
        );

    \I__4032\ : Odrv4
    port map (
            O => \N__25886\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__25883\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__4030\ : InMux
    port map (
            O => \N__25878\,
            I => \N__25875\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__25875\,
            I => \N__25871\
        );

    \I__4028\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25868\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__25871\,
            I => \N__25861\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__25868\,
            I => \N__25861\
        );

    \I__4025\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25858\
        );

    \I__4024\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25855\
        );

    \I__4023\ : Span4Mux_h
    port map (
            O => \N__25861\,
            I => \N__25850\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25850\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25847\
        );

    \I__4020\ : Odrv4
    port map (
            O => \N__25850\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__25847\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__4018\ : InMux
    port map (
            O => \N__25842\,
            I => \N__25836\
        );

    \I__4017\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25836\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__25836\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__4015\ : InMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__25830\,
            I => \N__25827\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__25827\,
            I => \N__25823\
        );

    \I__4012\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25820\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__25823\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__25820\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__25815\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\
        );

    \I__4008\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25806\
        );

    \I__4007\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25806\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__25806\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__4005\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25797\
        );

    \I__4004\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25797\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__25797\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__4002\ : InMux
    port map (
            O => \N__25794\,
            I => \N__25791\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__25791\,
            I => \N__25788\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__25788\,
            I => \N__25783\
        );

    \I__3999\ : InMux
    port map (
            O => \N__25787\,
            I => \N__25780\
        );

    \I__3998\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25777\
        );

    \I__3997\ : Span4Mux_v
    port map (
            O => \N__25783\,
            I => \N__25772\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__25780\,
            I => \N__25772\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__25777\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__25772\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__25767\,
            I => \N__25763\
        );

    \I__3992\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25758\
        );

    \I__3991\ : InMux
    port map (
            O => \N__25763\,
            I => \N__25758\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__25758\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__3989\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25749\
        );

    \I__3988\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25749\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__25749\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__25746\,
            I => \N__25742\
        );

    \I__3985\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25739\
        );

    \I__3984\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25736\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__25739\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__25736\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__3981\ : InMux
    port map (
            O => \N__25731\,
            I => \N__25727\
        );

    \I__3980\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25724\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__25727\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__25724\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__3977\ : InMux
    port map (
            O => \N__25719\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__3976\ : InMux
    port map (
            O => \N__25716\,
            I => \N__25713\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__25713\,
            I => \N__25709\
        );

    \I__3974\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25706\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__25709\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__25706\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__3971\ : CascadeMux
    port map (
            O => \N__25701\,
            I => \N__25696\
        );

    \I__3970\ : InMux
    port map (
            O => \N__25700\,
            I => \N__25693\
        );

    \I__3969\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25690\
        );

    \I__3968\ : InMux
    port map (
            O => \N__25696\,
            I => \N__25687\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__25693\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__25690\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__25687\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__3964\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__25677\,
            I => \N__25674\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__25674\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__3961\ : InMux
    port map (
            O => \N__25671\,
            I => \N__25665\
        );

    \I__3960\ : InMux
    port map (
            O => \N__25670\,
            I => \N__25665\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__25665\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__3957\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25653\
        );

    \I__3956\ : InMux
    port map (
            O => \N__25658\,
            I => \N__25653\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__25653\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__3954\ : InMux
    port map (
            O => \N__25650\,
            I => \N__25646\
        );

    \I__3953\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25643\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__25646\,
            I => \N__25640\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__25643\,
            I => \N__25637\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__25640\,
            I => \N__25634\
        );

    \I__3949\ : Span4Mux_h
    port map (
            O => \N__25637\,
            I => \N__25631\
        );

    \I__3948\ : Span4Mux_h
    port map (
            O => \N__25634\,
            I => \N__25628\
        );

    \I__3947\ : Span4Mux_h
    port map (
            O => \N__25631\,
            I => \N__25625\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__25628\,
            I => \N__25622\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__25625\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__25622\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__3943\ : InMux
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__25614\,
            I => \N__25611\
        );

    \I__3941\ : Span4Mux_v
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__3940\ : Sp12to4
    port map (
            O => \N__25608\,
            I => \N__25605\
        );

    \I__3939\ : Odrv12
    port map (
            O => \N__25605\,
            I => \pwm_generator_inst.O_12\
        );

    \I__3938\ : InMux
    port map (
            O => \N__25602\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__3937\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__25596\,
            I => \N__25593\
        );

    \I__3935\ : Span4Mux_v
    port map (
            O => \N__25593\,
            I => \N__25590\
        );

    \I__3934\ : Sp12to4
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__3933\ : Odrv12
    port map (
            O => \N__25587\,
            I => \pwm_generator_inst.O_13\
        );

    \I__3932\ : InMux
    port map (
            O => \N__25584\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__3931\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25578\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__3929\ : Sp12to4
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__3928\ : Span12Mux_s6_v
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__3927\ : Odrv12
    port map (
            O => \N__25569\,
            I => \pwm_generator_inst.O_14\
        );

    \I__3926\ : InMux
    port map (
            O => \N__25566\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__3925\ : InMux
    port map (
            O => \N__25563\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__3924\ : InMux
    port map (
            O => \N__25560\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__3923\ : InMux
    port map (
            O => \N__25557\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__3922\ : InMux
    port map (
            O => \N__25554\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__3921\ : InMux
    port map (
            O => \N__25551\,
            I => \bfn_9_27_0_\
        );

    \I__3920\ : CEMux
    port map (
            O => \N__25548\,
            I => \N__25543\
        );

    \I__3919\ : CEMux
    port map (
            O => \N__25547\,
            I => \N__25540\
        );

    \I__3918\ : CEMux
    port map (
            O => \N__25546\,
            I => \N__25537\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__25543\,
            I => \N__25533\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__25540\,
            I => \N__25530\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__25537\,
            I => \N__25527\
        );

    \I__3914\ : CEMux
    port map (
            O => \N__25536\,
            I => \N__25524\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__25533\,
            I => \N__25521\
        );

    \I__3912\ : Span4Mux_h
    port map (
            O => \N__25530\,
            I => \N__25518\
        );

    \I__3911\ : Span4Mux_h
    port map (
            O => \N__25527\,
            I => \N__25515\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__25524\,
            I => \N__25512\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__25521\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__25518\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__25515\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__3906\ : Odrv12
    port map (
            O => \N__25512\,
            I => \delay_measurement_inst.delay_hc_timer.N_199_i\
        );

    \I__3905\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25500\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__25500\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__3903\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25493\
        );

    \I__3902\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25490\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__25493\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25490\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25482\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__25482\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__3897\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__25476\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__25473\,
            I => \N__25468\
        );

    \I__3894\ : InMux
    port map (
            O => \N__25472\,
            I => \N__25465\
        );

    \I__3893\ : InMux
    port map (
            O => \N__25471\,
            I => \N__25462\
        );

    \I__3892\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25459\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25465\,
            I => \current_shift_inst.N_1288_i\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__25462\,
            I => \current_shift_inst.N_1288_i\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__25459\,
            I => \current_shift_inst.N_1288_i\
        );

    \I__3888\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__25449\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25446\,
            I => \N__25443\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__25443\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3883\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25431\
        );

    \I__3882\ : InMux
    port map (
            O => \N__25436\,
            I => \N__25431\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__25428\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__3879\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25419\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25419\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25419\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__3876\ : InMux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__3874\ : Span4Mux_h
    port map (
            O => \N__25410\,
            I => \N__25406\
        );

    \I__3873\ : InMux
    port map (
            O => \N__25409\,
            I => \N__25403\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__25406\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__25403\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__25398\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\
        );

    \I__3869\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25390\
        );

    \I__3868\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25385\
        );

    \I__3867\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25385\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__25390\,
            I => \N__25381\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__25385\,
            I => \N__25378\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25375\
        );

    \I__3863\ : Span4Mux_v
    port map (
            O => \N__25381\,
            I => \N__25370\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__25378\,
            I => \N__25370\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__25375\,
            I => \N__25367\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__25370\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__25367\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25359\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__3856\ : Span12Mux_v
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3855\ : Odrv12
    port map (
            O => \N__25353\,
            I => il_min_comp1_c
        );

    \I__3854\ : InMux
    port map (
            O => \N__25350\,
            I => \N__25338\
        );

    \I__3853\ : InMux
    port map (
            O => \N__25349\,
            I => \N__25338\
        );

    \I__3852\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25338\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25338\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__25338\,
            I => \N__25309\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25337\,
            I => \N__25300\
        );

    \I__3848\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25300\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25335\,
            I => \N__25300\
        );

    \I__3846\ : InMux
    port map (
            O => \N__25334\,
            I => \N__25300\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25295\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25295\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25286\
        );

    \I__3842\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25286\
        );

    \I__3841\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25286\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25328\,
            I => \N__25286\
        );

    \I__3839\ : InMux
    port map (
            O => \N__25327\,
            I => \N__25277\
        );

    \I__3838\ : InMux
    port map (
            O => \N__25326\,
            I => \N__25277\
        );

    \I__3837\ : InMux
    port map (
            O => \N__25325\,
            I => \N__25277\
        );

    \I__3836\ : InMux
    port map (
            O => \N__25324\,
            I => \N__25277\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25323\,
            I => \N__25268\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25322\,
            I => \N__25268\
        );

    \I__3833\ : InMux
    port map (
            O => \N__25321\,
            I => \N__25268\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25268\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25259\
        );

    \I__3830\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25259\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25259\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25316\,
            I => \N__25259\
        );

    \I__3827\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25250\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25250\
        );

    \I__3825\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25250\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25250\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__25309\,
            I => \N__25247\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__25300\,
            I => \N__25244\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__25295\,
            I => \N__25241\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25234\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25277\,
            I => \N__25234\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25268\,
            I => \N__25234\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__25259\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25250\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__25247\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__25244\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3813\ : Odrv4
    port map (
            O => \N__25241\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__25234\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__3811\ : CEMux
    port map (
            O => \N__25221\,
            I => \N__25214\
        );

    \I__3810\ : CEMux
    port map (
            O => \N__25220\,
            I => \N__25211\
        );

    \I__3809\ : CEMux
    port map (
            O => \N__25219\,
            I => \N__25208\
        );

    \I__3808\ : CEMux
    port map (
            O => \N__25218\,
            I => \N__25205\
        );

    \I__3807\ : CEMux
    port map (
            O => \N__25217\,
            I => \N__25202\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__25214\,
            I => \N__25199\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25211\,
            I => \N__25196\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__25208\,
            I => \N__25193\
        );

    \I__3803\ : LocalMux
    port map (
            O => \N__25205\,
            I => \N__25190\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__25202\,
            I => \N__25187\
        );

    \I__3801\ : Span4Mux_h
    port map (
            O => \N__25199\,
            I => \N__25184\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__25196\,
            I => \N__25181\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__25193\,
            I => \N__25176\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__25190\,
            I => \N__25176\
        );

    \I__3797\ : Span4Mux_h
    port map (
            O => \N__25187\,
            I => \N__25173\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__25184\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__3795\ : Odrv4
    port map (
            O => \N__25181\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__25176\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__25173\,
            I => \delay_measurement_inst.delay_hc_timer.N_198_i\
        );

    \I__3792\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25160\
        );

    \I__3791\ : InMux
    port map (
            O => \N__25163\,
            I => \N__25156\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__25160\,
            I => \N__25153\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25150\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25156\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__25153\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25150\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__3785\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25140\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25140\,
            I => \N__25136\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25139\,
            I => \N__25133\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__25136\,
            I => \N__25128\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__25133\,
            I => \N__25128\
        );

    \I__3780\ : Span4Mux_v
    port map (
            O => \N__25128\,
            I => \N__25123\
        );

    \I__3779\ : InMux
    port map (
            O => \N__25127\,
            I => \N__25120\
        );

    \I__3778\ : InMux
    port map (
            O => \N__25126\,
            I => \N__25117\
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__25123\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__25120\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__25117\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__3774\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25104\
        );

    \I__3773\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25104\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25104\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25097\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25094\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25090\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25094\,
            I => \N__25087\
        );

    \I__3767\ : InMux
    port map (
            O => \N__25093\,
            I => \N__25084\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__25090\,
            I => \N__25081\
        );

    \I__3765\ : Span4Mux_h
    port map (
            O => \N__25087\,
            I => \N__25078\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__25084\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__3763\ : Odrv4
    port map (
            O => \N__25081\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__25078\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__25071\,
            I => \N__25065\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25070\,
            I => \N__25062\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25059\
        );

    \I__3758\ : InMux
    port map (
            O => \N__25068\,
            I => \N__25056\
        );

    \I__3757\ : InMux
    port map (
            O => \N__25065\,
            I => \N__25053\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__25062\,
            I => \N__25050\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__25059\,
            I => \N__25047\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25042\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__25053\,
            I => \N__25042\
        );

    \I__3752\ : Span4Mux_h
    port map (
            O => \N__25050\,
            I => \N__25039\
        );

    \I__3751\ : Span4Mux_h
    port map (
            O => \N__25047\,
            I => \N__25034\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__25042\,
            I => \N__25034\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__25039\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__25034\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__25029\,
            I => \N__25026\
        );

    \I__3746\ : InMux
    port map (
            O => \N__25026\,
            I => \N__25020\
        );

    \I__3745\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25020\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25020\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25017\,
            I => \N__25012\
        );

    \I__3742\ : InMux
    port map (
            O => \N__25016\,
            I => \N__25006\
        );

    \I__3741\ : InMux
    port map (
            O => \N__25015\,
            I => \N__25006\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__25012\,
            I => \N__25003\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25011\,
            I => \N__25000\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25006\,
            I => \N__24997\
        );

    \I__3737\ : Span4Mux_h
    port map (
            O => \N__25003\,
            I => \N__24992\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25000\,
            I => \N__24992\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__24997\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__24992\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__3733\ : InMux
    port map (
            O => \N__24987\,
            I => \N__24984\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__24984\,
            I => \N__24981\
        );

    \I__3731\ : Span4Mux_h
    port map (
            O => \N__24981\,
            I => \N__24977\
        );

    \I__3730\ : InMux
    port map (
            O => \N__24980\,
            I => \N__24974\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__24977\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__24974\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__3727\ : InMux
    port map (
            O => \N__24969\,
            I => \N__24966\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__24966\,
            I => \N__24962\
        );

    \I__3725\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24958\
        );

    \I__3724\ : Span4Mux_v
    port map (
            O => \N__24962\,
            I => \N__24955\
        );

    \I__3723\ : InMux
    port map (
            O => \N__24961\,
            I => \N__24952\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__24958\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__24955\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__24952\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__3719\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24941\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__24944\,
            I => \N__24936\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__24941\,
            I => \N__24933\
        );

    \I__3716\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24930\
        );

    \I__3715\ : InMux
    port map (
            O => \N__24939\,
            I => \N__24927\
        );

    \I__3714\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24924\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__24933\,
            I => \N__24921\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__24930\,
            I => \N__24916\
        );

    \I__3711\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24916\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24913\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__24921\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__24916\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__24913\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__3706\ : InMux
    port map (
            O => \N__24906\,
            I => \N__24902\
        );

    \I__3705\ : InMux
    port map (
            O => \N__24905\,
            I => \N__24898\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__24902\,
            I => \N__24895\
        );

    \I__3703\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24892\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__24898\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__3701\ : Odrv12
    port map (
            O => \N__24895\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__24892\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__3699\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24880\
        );

    \I__3698\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24877\
        );

    \I__3697\ : InMux
    port map (
            O => \N__24883\,
            I => \N__24874\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__24880\,
            I => \N__24870\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__24877\,
            I => \N__24867\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__24874\,
            I => \N__24864\
        );

    \I__3693\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24861\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__24870\,
            I => \N__24856\
        );

    \I__3691\ : Span4Mux_v
    port map (
            O => \N__24867\,
            I => \N__24856\
        );

    \I__3690\ : Span4Mux_h
    port map (
            O => \N__24864\,
            I => \N__24851\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__24861\,
            I => \N__24851\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__24856\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__24851\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__3686\ : InMux
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__24843\,
            I => \N__24837\
        );

    \I__3684\ : InMux
    port map (
            O => \N__24842\,
            I => \N__24834\
        );

    \I__3683\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24831\
        );

    \I__3682\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24828\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__24837\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__24834\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__24831\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__24828\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__3677\ : InMux
    port map (
            O => \N__24819\,
            I => \N__24815\
        );

    \I__3676\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24811\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24808\
        );

    \I__3674\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24805\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__24811\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__24808\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__24805\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__3670\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24794\
        );

    \I__3669\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24790\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__24794\,
            I => \N__24787\
        );

    \I__3667\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24784\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__24790\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__3665\ : Odrv12
    port map (
            O => \N__24787\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__24784\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__3663\ : InMux
    port map (
            O => \N__24777\,
            I => \N__24773\
        );

    \I__3662\ : InMux
    port map (
            O => \N__24776\,
            I => \N__24769\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24765\
        );

    \I__3660\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24762\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__24769\,
            I => \N__24759\
        );

    \I__3658\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24756\
        );

    \I__3657\ : Span4Mux_h
    port map (
            O => \N__24765\,
            I => \N__24753\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24750\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__24759\,
            I => \N__24747\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__24756\,
            I => \N__24744\
        );

    \I__3653\ : Span4Mux_v
    port map (
            O => \N__24753\,
            I => \N__24741\
        );

    \I__3652\ : Span4Mux_h
    port map (
            O => \N__24750\,
            I => \N__24738\
        );

    \I__3651\ : Span4Mux_v
    port map (
            O => \N__24747\,
            I => \N__24733\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__24744\,
            I => \N__24733\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__24741\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__24738\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__24733\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__3646\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24723\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__24723\,
            I => \N__24719\
        );

    \I__3644\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24715\
        );

    \I__3643\ : Span4Mux_v
    port map (
            O => \N__24719\,
            I => \N__24712\
        );

    \I__3642\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24709\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__24715\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__24712\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__24709\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__3638\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24698\
        );

    \I__3637\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24693\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__24698\,
            I => \N__24690\
        );

    \I__3635\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24685\
        );

    \I__3634\ : InMux
    port map (
            O => \N__24696\,
            I => \N__24685\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24682\
        );

    \I__3632\ : Span4Mux_h
    port map (
            O => \N__24690\,
            I => \N__24679\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__24685\,
            I => \N__24676\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__24682\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__24679\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__24676\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__3627\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24665\
        );

    \I__3626\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24662\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__24665\,
            I => \N__24657\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__24662\,
            I => \N__24654\
        );

    \I__3623\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24649\
        );

    \I__3622\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24649\
        );

    \I__3621\ : Span4Mux_v
    port map (
            O => \N__24657\,
            I => \N__24642\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__24654\,
            I => \N__24642\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__24649\,
            I => \N__24642\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__24642\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__3617\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24634\
        );

    \I__3616\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24631\
        );

    \I__3615\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24628\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__24634\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__24631\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__24628\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__3611\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24617\
        );

    \I__3610\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24614\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__24617\,
            I => \N__24609\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__24614\,
            I => \N__24606\
        );

    \I__3607\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24601\
        );

    \I__3606\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24601\
        );

    \I__3605\ : Span4Mux_v
    port map (
            O => \N__24609\,
            I => \N__24598\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__24606\,
            I => \N__24593\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__24601\,
            I => \N__24593\
        );

    \I__3602\ : Span4Mux_v
    port map (
            O => \N__24598\,
            I => \N__24590\
        );

    \I__3601\ : Span4Mux_v
    port map (
            O => \N__24593\,
            I => \N__24587\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__24590\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__24587\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__3598\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24578\
        );

    \I__3597\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24574\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__24578\,
            I => \N__24571\
        );

    \I__3595\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24568\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__24574\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__24571\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__24568\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__3591\ : InMux
    port map (
            O => \N__24561\,
            I => \N__24557\
        );

    \I__3590\ : InMux
    port map (
            O => \N__24560\,
            I => \N__24553\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__24557\,
            I => \N__24550\
        );

    \I__3588\ : InMux
    port map (
            O => \N__24556\,
            I => \N__24547\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__24553\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__3586\ : Odrv4
    port map (
            O => \N__24550\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__24547\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__3584\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__24537\,
            I => \N__24533\
        );

    \I__3582\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24530\
        );

    \I__3581\ : Span4Mux_v
    port map (
            O => \N__24533\,
            I => \N__24526\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24523\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__24529\,
            I => \N__24519\
        );

    \I__3578\ : Span4Mux_h
    port map (
            O => \N__24526\,
            I => \N__24516\
        );

    \I__3577\ : Span4Mux_h
    port map (
            O => \N__24523\,
            I => \N__24513\
        );

    \I__3576\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24508\
        );

    \I__3575\ : InMux
    port map (
            O => \N__24519\,
            I => \N__24508\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__24516\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__3573\ : Odrv4
    port map (
            O => \N__24513\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__24508\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__24501\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__3569\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24489\
        );

    \I__3568\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24489\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__24489\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__3566\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24480\
        );

    \I__3565\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24480\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__24480\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__3563\ : IoInMux
    port map (
            O => \N__24477\,
            I => \N__24474\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__24474\,
            I => \GB_BUFFER_clock_output_0_THRU_CO\
        );

    \I__3561\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__24468\,
            I => \N__24465\
        );

    \I__3559\ : Glb2LocalMux
    port map (
            O => \N__24465\,
            I => \N__24462\
        );

    \I__3558\ : GlobalMux
    port map (
            O => \N__24462\,
            I => clk_12mhz
        );

    \I__3557\ : IoInMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24453\
        );

    \I__3555\ : Span4Mux_s0_v
    port map (
            O => \N__24453\,
            I => \N__24450\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__24450\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__3553\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24444\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__24444\,
            I => \N__24441\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__24441\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24438\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__3549\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24432\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__24432\,
            I => \N__24429\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__24429\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24426\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__24420\,
            I => \N__24417\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__24417\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24414\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__3541\ : InMux
    port map (
            O => \N__24411\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__3540\ : InMux
    port map (
            O => \N__24408\,
            I => \N__24405\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__24405\,
            I => \N__24401\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24404\,
            I => \N__24398\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__24401\,
            I => \current_shift_inst.control_input_31\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__24398\,
            I => \current_shift_inst.control_input_31\
        );

    \I__3535\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__24390\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__3531\ : Span4Mux_h
    port map (
            O => \N__24381\,
            I => \N__24377\
        );

    \I__3530\ : InMux
    port map (
            O => \N__24380\,
            I => \N__24374\
        );

    \I__3529\ : Span4Mux_v
    port map (
            O => \N__24377\,
            I => \N__24371\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__24374\,
            I => \N__24368\
        );

    \I__3527\ : Span4Mux_h
    port map (
            O => \N__24371\,
            I => \N__24365\
        );

    \I__3526\ : Odrv12
    port map (
            O => \N__24368\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__24365\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__3524\ : IoInMux
    port map (
            O => \N__24360\,
            I => \N__24357\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__3522\ : Span12Mux_s7_v
    port map (
            O => \N__24354\,
            I => \N__24351\
        );

    \I__3521\ : Odrv12
    port map (
            O => \N__24351\,
            I => s4_phy_c
        );

    \I__3520\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__24342\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24339\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24333\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24330\
        );

    \I__3514\ : Odrv4
    port map (
            O => \N__24330\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24327\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__24318\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24315\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24309\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__24309\,
            I => \N__24306\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__24306\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__3505\ : InMux
    port map (
            O => \N__24303\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__3504\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__3502\ : Odrv12
    port map (
            O => \N__24294\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__3501\ : InMux
    port map (
            O => \N__24291\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__3500\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__24285\,
            I => \N__24282\
        );

    \I__3498\ : Odrv12
    port map (
            O => \N__24282\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__3497\ : InMux
    port map (
            O => \N__24279\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24276\,
            I => \N__24273\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24270\
        );

    \I__3494\ : Odrv12
    port map (
            O => \N__24270\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24267\,
            I => \bfn_8_16_0_\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24261\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__24261\,
            I => \N__24258\
        );

    \I__3490\ : Odrv12
    port map (
            O => \N__24258\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__3489\ : InMux
    port map (
            O => \N__24255\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__24252\,
            I => \N__24248\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__24251\,
            I => \N__24245\
        );

    \I__3486\ : InMux
    port map (
            O => \N__24248\,
            I => \N__24241\
        );

    \I__3485\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24238\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24235\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__24241\,
            I => \N__24232\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__24238\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24235\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__24232\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24225\,
            I => \bfn_8_14_0_\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__24222\,
            I => \N__24218\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__24221\,
            I => \N__24215\
        );

    \I__3476\ : InMux
    port map (
            O => \N__24218\,
            I => \N__24211\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24215\,
            I => \N__24208\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24205\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24211\,
            I => \N__24202\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24208\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24205\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__24202\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__3469\ : InMux
    port map (
            O => \N__24195\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__24192\,
            I => \N__24189\
        );

    \I__3467\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24184\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24181\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24178\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__24184\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24181\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__24178\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24171\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__24168\,
            I => \N__24165\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24160\
        );

    \I__3458\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24157\
        );

    \I__3457\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24154\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__24160\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__24157\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24154\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24147\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24140\
        );

    \I__3451\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24137\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__24140\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__24137\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__3448\ : InMux
    port map (
            O => \N__24132\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__3447\ : InMux
    port map (
            O => \N__24129\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__3446\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24122\
        );

    \I__3445\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24119\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__24122\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24119\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__3442\ : InMux
    port map (
            O => \N__24114\,
            I => \N__24111\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__24111\,
            I => \N__24108\
        );

    \I__3440\ : Odrv12
    port map (
            O => \N__24108\,
            I => \current_shift_inst.control_input_18\
        );

    \I__3439\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24102\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__24102\,
            I => \N__24099\
        );

    \I__3437\ : Odrv12
    port map (
            O => \N__24099\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__3436\ : InMux
    port map (
            O => \N__24096\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24088\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24083\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24091\,
            I => \N__24083\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__24088\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24083\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__3430\ : InMux
    port map (
            O => \N__24078\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__24075\,
            I => \N__24071\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__24074\,
            I => \N__24068\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24071\,
            I => \N__24064\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24061\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24067\,
            I => \N__24058\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24064\,
            I => \N__24055\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24061\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24058\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__24055\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24048\,
            I => \bfn_8_13_0_\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__24045\,
            I => \N__24041\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__24044\,
            I => \N__24038\
        );

    \I__3417\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24034\
        );

    \I__3416\ : InMux
    port map (
            O => \N__24038\,
            I => \N__24031\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24028\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24034\,
            I => \N__24025\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__24031\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__24028\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__3411\ : Odrv4
    port map (
            O => \N__24025\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__3410\ : InMux
    port map (
            O => \N__24018\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24010\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24014\,
            I => \N__24005\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24005\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24010\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__24005\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__3404\ : InMux
    port map (
            O => \N__24000\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__3402\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23989\
        );

    \I__3401\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23986\
        );

    \I__3400\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23983\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__23989\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__23986\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__23983\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__3396\ : InMux
    port map (
            O => \N__23976\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__23973\,
            I => \N__23968\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__23972\,
            I => \N__23965\
        );

    \I__3393\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23962\
        );

    \I__3392\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23957\
        );

    \I__3391\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23957\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__23962\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__23957\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__3388\ : InMux
    port map (
            O => \N__23952\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__23949\,
            I => \N__23946\
        );

    \I__3386\ : InMux
    port map (
            O => \N__23946\,
            I => \N__23941\
        );

    \I__3385\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23938\
        );

    \I__3384\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23935\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__23941\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__23938\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__23935\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__3380\ : InMux
    port map (
            O => \N__23928\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__3379\ : InMux
    port map (
            O => \N__23925\,
            I => \N__23920\
        );

    \I__3378\ : InMux
    port map (
            O => \N__23924\,
            I => \N__23915\
        );

    \I__3377\ : InMux
    port map (
            O => \N__23923\,
            I => \N__23915\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__23920\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__23915\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__3374\ : InMux
    port map (
            O => \N__23910\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__3373\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23902\
        );

    \I__3372\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23897\
        );

    \I__3371\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23897\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__23902\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__23897\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__3368\ : InMux
    port map (
            O => \N__23892\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__3367\ : InMux
    port map (
            O => \N__23889\,
            I => \N__23884\
        );

    \I__3366\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23879\
        );

    \I__3365\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23879\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__23884\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__23879\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__3362\ : InMux
    port map (
            O => \N__23874\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__23871\,
            I => \N__23867\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__23870\,
            I => \N__23864\
        );

    \I__3359\ : InMux
    port map (
            O => \N__23867\,
            I => \N__23860\
        );

    \I__3358\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23857\
        );

    \I__3357\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23854\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23851\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__23857\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__23854\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__23851\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__3352\ : InMux
    port map (
            O => \N__23844\,
            I => \bfn_8_12_0_\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__23841\,
            I => \N__23837\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__23840\,
            I => \N__23834\
        );

    \I__3349\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23830\
        );

    \I__3348\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23827\
        );

    \I__3347\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23824\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23821\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__23827\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__23824\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__23821\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__3342\ : InMux
    port map (
            O => \N__23814\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__3341\ : InMux
    port map (
            O => \N__23811\,
            I => \N__23806\
        );

    \I__3340\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23801\
        );

    \I__3339\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23801\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__23806\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__23801\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__3336\ : InMux
    port map (
            O => \N__23796\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__23793\,
            I => \N__23790\
        );

    \I__3334\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23785\
        );

    \I__3333\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23782\
        );

    \I__3332\ : InMux
    port map (
            O => \N__23788\,
            I => \N__23779\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__23785\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__23782\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__23779\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__3328\ : InMux
    port map (
            O => \N__23772\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__23769\,
            I => \N__23764\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__23768\,
            I => \N__23761\
        );

    \I__3325\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23758\
        );

    \I__3324\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23753\
        );

    \I__3323\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23753\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__23758\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__23753\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__3320\ : InMux
    port map (
            O => \N__23748\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__3318\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23737\
        );

    \I__3317\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23734\
        );

    \I__3316\ : InMux
    port map (
            O => \N__23740\,
            I => \N__23731\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__23737\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__23734\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__23731\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__3312\ : InMux
    port map (
            O => \N__23724\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__3311\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23716\
        );

    \I__3310\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23711\
        );

    \I__3309\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23711\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__23716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__23711\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__3306\ : InMux
    port map (
            O => \N__23706\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__23703\,
            I => \N__23699\
        );

    \I__3304\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23695\
        );

    \I__3303\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23692\
        );

    \I__3302\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23689\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__23695\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__23692\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__23689\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__3298\ : InMux
    port map (
            O => \N__23682\,
            I => \bfn_8_11_0_\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__23679\,
            I => \N__23675\
        );

    \I__3296\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23671\
        );

    \I__3295\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23668\
        );

    \I__3294\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23665\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__23671\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__23668\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__23665\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__3290\ : InMux
    port map (
            O => \N__23658\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__3289\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23650\
        );

    \I__3288\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23645\
        );

    \I__3287\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23645\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__23650\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__23645\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__3284\ : InMux
    port map (
            O => \N__23640\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__23637\,
            I => \N__23634\
        );

    \I__3282\ : InMux
    port map (
            O => \N__23634\,
            I => \N__23629\
        );

    \I__3281\ : InMux
    port map (
            O => \N__23633\,
            I => \N__23626\
        );

    \I__3280\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23623\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__23629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__23626\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__23623\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__3276\ : InMux
    port map (
            O => \N__23616\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__23613\,
            I => \N__23608\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__23612\,
            I => \N__23605\
        );

    \I__3273\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23602\
        );

    \I__3272\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23597\
        );

    \I__3271\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23597\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__23602\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__23597\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__3268\ : InMux
    port map (
            O => \N__23592\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__23589\,
            I => \N__23586\
        );

    \I__3266\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23581\
        );

    \I__3265\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23578\
        );

    \I__3264\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23575\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__23581\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__23578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__23575\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__3260\ : InMux
    port map (
            O => \N__23568\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__3259\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23560\
        );

    \I__3258\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23555\
        );

    \I__3257\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23555\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__23560\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__23555\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__3254\ : InMux
    port map (
            O => \N__23550\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__3253\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23544\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__23544\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__3251\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23538\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__23538\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\
        );

    \I__3249\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23532\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__23532\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\
        );

    \I__3247\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23526\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__23526\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__3245\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23519\
        );

    \I__3244\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23516\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__23519\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__23516\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__3241\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23505\
        );

    \I__3240\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23505\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__23505\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__23502\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\
        );

    \I__3237\ : InMux
    port map (
            O => \N__23499\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__3236\ : InMux
    port map (
            O => \N__23496\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__3235\ : InMux
    port map (
            O => \N__23493\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23490\,
            I => \bfn_7_28_0_\
        );

    \I__3233\ : InMux
    port map (
            O => \N__23487\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__3232\ : InMux
    port map (
            O => \N__23484\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23481\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__3230\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23475\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23472\
        );

    \I__3228\ : Odrv12
    port map (
            O => \N__23472\,
            I => il_max_comp1_c
        );

    \I__3227\ : InMux
    port map (
            O => \N__23469\,
            I => \N__23466\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__23466\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__3225\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23460\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__23460\,
            I => \N__23457\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__23457\,
            I => \N__23454\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__23454\,
            I => \N__23451\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__23451\,
            I => \pwm_generator_inst.O_5\
        );

    \I__3220\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23445\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__23445\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23439\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__23439\,
            I => \N__23436\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__23436\,
            I => \N__23433\
        );

    \I__3215\ : Span4Mux_h
    port map (
            O => \N__23433\,
            I => \N__23430\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__23430\,
            I => \pwm_generator_inst.O_6\
        );

    \I__3213\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23424\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23424\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23418\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23415\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__23415\,
            I => \N__23412\
        );

    \I__3208\ : Span4Mux_h
    port map (
            O => \N__23412\,
            I => \N__23409\
        );

    \I__3207\ : Odrv4
    port map (
            O => \N__23409\,
            I => \pwm_generator_inst.O_7\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23403\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__23403\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__3204\ : InMux
    port map (
            O => \N__23400\,
            I => \N__23397\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__23397\,
            I => \N__23394\
        );

    \I__3202\ : Span4Mux_v
    port map (
            O => \N__23394\,
            I => \N__23391\
        );

    \I__3201\ : Span4Mux_h
    port map (
            O => \N__23391\,
            I => \N__23388\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__23388\,
            I => \pwm_generator_inst.O_8\
        );

    \I__3199\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__23382\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__3197\ : InMux
    port map (
            O => \N__23379\,
            I => \N__23376\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23376\,
            I => \N__23373\
        );

    \I__3195\ : Span12Mux_s6_v
    port map (
            O => \N__23373\,
            I => \N__23370\
        );

    \I__3194\ : Odrv12
    port map (
            O => \N__23370\,
            I => \pwm_generator_inst.O_9\
        );

    \I__3193\ : InMux
    port map (
            O => \N__23367\,
            I => \N__23364\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23364\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__3191\ : InMux
    port map (
            O => \N__23361\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__3190\ : InMux
    port map (
            O => \N__23358\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__3189\ : InMux
    port map (
            O => \N__23355\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23349\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23346\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__23346\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__3185\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23340\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__23340\,
            I => \N__23337\
        );

    \I__3183\ : Span4Mux_v
    port map (
            O => \N__23337\,
            I => \N__23334\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__23334\,
            I => \N__23331\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__23331\,
            I => \pwm_generator_inst.O_0\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__23328\,
            I => \N__23325\
        );

    \I__3179\ : InMux
    port map (
            O => \N__23325\,
            I => \N__23322\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__23322\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__3177\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23316\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__23316\,
            I => \N__23313\
        );

    \I__3175\ : Span12Mux_s7_v
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__3174\ : Odrv12
    port map (
            O => \N__23310\,
            I => \pwm_generator_inst.O_1\
        );

    \I__3173\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23304\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__23304\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__3171\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23298\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__23298\,
            I => \N__23295\
        );

    \I__3169\ : Span4Mux_h
    port map (
            O => \N__23295\,
            I => \N__23292\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__23292\,
            I => \N__23289\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__23289\,
            I => \pwm_generator_inst.O_2\
        );

    \I__3166\ : InMux
    port map (
            O => \N__23286\,
            I => \N__23283\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__23283\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23277\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23277\,
            I => \N__23274\
        );

    \I__3162\ : Span4Mux_h
    port map (
            O => \N__23274\,
            I => \N__23271\
        );

    \I__3161\ : Span4Mux_h
    port map (
            O => \N__23271\,
            I => \N__23268\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__23268\,
            I => \pwm_generator_inst.O_3\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23262\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__3157\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23256\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__3155\ : Span4Mux_h
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__23250\,
            I => \N__23247\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__23247\,
            I => \pwm_generator_inst.O_4\
        );

    \I__3152\ : InMux
    port map (
            O => \N__23244\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23241\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23238\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__3149\ : InMux
    port map (
            O => \N__23235\,
            I => \bfn_7_13_0_\
        );

    \I__3148\ : InMux
    port map (
            O => \N__23232\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23229\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23226\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23223\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23220\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23217\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3142\ : InMux
    port map (
            O => \N__23214\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23211\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23208\,
            I => \bfn_7_12_0_\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23205\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__3138\ : InMux
    port map (
            O => \N__23202\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__3137\ : InMux
    port map (
            O => \N__23199\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__3136\ : InMux
    port map (
            O => \N__23196\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3135\ : InMux
    port map (
            O => \N__23193\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23190\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23187\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23184\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23181\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3130\ : InMux
    port map (
            O => \N__23178\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3129\ : InMux
    port map (
            O => \N__23175\,
            I => \bfn_7_11_0_\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23172\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23169\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23166\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__3125\ : InMux
    port map (
            O => \N__23163\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__3124\ : InMux
    port map (
            O => \N__23160\,
            I => \N__23128\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23128\
        );

    \I__3122\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23128\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23128\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23128\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23155\,
            I => \N__23128\
        );

    \I__3118\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23128\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23128\
        );

    \I__3116\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23111\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23111\
        );

    \I__3114\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23111\
        );

    \I__3113\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23111\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23111\
        );

    \I__3111\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23111\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23111\
        );

    \I__3109\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23111\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23107\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23111\,
            I => \N__23104\
        );

    \I__3106\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23101\
        );

    \I__3105\ : Span4Mux_v
    port map (
            O => \N__23107\,
            I => \N__23098\
        );

    \I__3104\ : Span4Mux_v
    port map (
            O => \N__23104\,
            I => \N__23095\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23092\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__23098\,
            I => \N__23086\
        );

    \I__3101\ : Span4Mux_v
    port map (
            O => \N__23095\,
            I => \N__23086\
        );

    \I__3100\ : Span4Mux_s2_h
    port map (
            O => \N__23092\,
            I => \N__23083\
        );

    \I__3099\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23080\
        );

    \I__3098\ : Span4Mux_h
    port map (
            O => \N__23086\,
            I => \N__23077\
        );

    \I__3097\ : Span4Mux_v
    port map (
            O => \N__23083\,
            I => \N__23074\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__23080\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__23077\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__23074\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23063\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23060\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23063\,
            I => \N__23057\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__23060\,
            I => \N__23054\
        );

    \I__3089\ : Span12Mux_v
    port map (
            O => \N__23057\,
            I => \N__23051\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__23054\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__3087\ : Odrv12
    port map (
            O => \N__23051\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23043\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__23043\,
            I => \N__23040\
        );

    \I__3084\ : Odrv12
    port map (
            O => \N__23040\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__23037\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\
        );

    \I__3082\ : InMux
    port map (
            O => \N__23034\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3081\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__23024\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23027\,
            I => \N__23021\
        );

    \I__3078\ : Span4Mux_s1_h
    port map (
            O => \N__23024\,
            I => \N__23018\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23021\,
            I => \N__23015\
        );

    \I__3076\ : Span4Mux_h
    port map (
            O => \N__23018\,
            I => \N__23012\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__23015\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__23012\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23007\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__3072\ : InMux
    port map (
            O => \N__23004\,
            I => \N__23000\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22997\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22994\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22991\
        );

    \I__3068\ : Span4Mux_s1_h
    port map (
            O => \N__22994\,
            I => \N__22988\
        );

    \I__3067\ : Span4Mux_h
    port map (
            O => \N__22991\,
            I => \N__22983\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__22988\,
            I => \N__22983\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__22983\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__3064\ : InMux
    port map (
            O => \N__22980\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__3063\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22974\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__22974\,
            I => \N__22970\
        );

    \I__3061\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22967\
        );

    \I__3060\ : Span12Mux_s5_h
    port map (
            O => \N__22970\,
            I => \N__22964\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__22967\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__3058\ : Odrv12
    port map (
            O => \N__22964\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__3057\ : InMux
    port map (
            O => \N__22959\,
            I => \bfn_5_16_0_\
        );

    \I__3056\ : InMux
    port map (
            O => \N__22956\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__3055\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22950\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__22950\,
            I => \N__22946\
        );

    \I__3053\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22943\
        );

    \I__3052\ : Span4Mux_s1_h
    port map (
            O => \N__22946\,
            I => \N__22940\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__22943\,
            I => \N__22937\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__22940\,
            I => \N__22934\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__22937\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__22934\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__3047\ : InMux
    port map (
            O => \N__22929\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__3046\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22923\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__22923\,
            I => \N__22919\
        );

    \I__3044\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22916\
        );

    \I__3043\ : Span4Mux_s1_h
    port map (
            O => \N__22919\,
            I => \N__22913\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22910\
        );

    \I__3041\ : Span4Mux_h
    port map (
            O => \N__22913\,
            I => \N__22907\
        );

    \I__3040\ : Odrv4
    port map (
            O => \N__22910\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__3039\ : Odrv4
    port map (
            O => \N__22907\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__3038\ : InMux
    port map (
            O => \N__22902\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__3037\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__22896\,
            I => \N__22893\
        );

    \I__3035\ : Span4Mux_s1_h
    port map (
            O => \N__22893\,
            I => \N__22889\
        );

    \I__3034\ : InMux
    port map (
            O => \N__22892\,
            I => \N__22886\
        );

    \I__3033\ : Span4Mux_h
    port map (
            O => \N__22889\,
            I => \N__22883\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__22886\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__3031\ : Odrv4
    port map (
            O => \N__22883\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__3030\ : InMux
    port map (
            O => \N__22878\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__3029\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22872\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__22872\,
            I => \N__22868\
        );

    \I__3027\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22865\
        );

    \I__3026\ : Span4Mux_s1_h
    port map (
            O => \N__22868\,
            I => \N__22862\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__22865\,
            I => \N__22859\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__22862\,
            I => \N__22856\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__22859\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3022\ : Odrv4
    port map (
            O => \N__22856\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__3021\ : InMux
    port map (
            O => \N__22851\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__3020\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__22842\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__3017\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__22836\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__3015\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22828\
        );

    \I__3014\ : InMux
    port map (
            O => \N__22832\,
            I => \N__22825\
        );

    \I__3013\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22822\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__22828\,
            I => \N__22819\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__22825\,
            I => \N__22816\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__22822\,
            I => \N__22812\
        );

    \I__3009\ : Span4Mux_v
    port map (
            O => \N__22819\,
            I => \N__22809\
        );

    \I__3008\ : Span4Mux_v
    port map (
            O => \N__22816\,
            I => \N__22806\
        );

    \I__3007\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22803\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__22812\,
            I => \N__22800\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__22809\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__22806\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__22803\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__22800\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__3001\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22787\
        );

    \I__3000\ : InMux
    port map (
            O => \N__22790\,
            I => \N__22783\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22780\
        );

    \I__2998\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22777\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__22783\,
            I => \N__22774\
        );

    \I__2996\ : Span4Mux_h
    port map (
            O => \N__22780\,
            I => \N__22768\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__22777\,
            I => \N__22768\
        );

    \I__2994\ : Span4Mux_h
    port map (
            O => \N__22774\,
            I => \N__22765\
        );

    \I__2993\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22762\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__22768\,
            I => \N__22759\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__22765\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__22762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__22759\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__22752\,
            I => \N__22748\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__22751\,
            I => \N__22745\
        );

    \I__2986\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22741\
        );

    \I__2985\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22738\
        );

    \I__2984\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22734\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__22741\,
            I => \N__22731\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__22738\,
            I => \N__22728\
        );

    \I__2981\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22725\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22722\
        );

    \I__2979\ : Span4Mux_h
    port map (
            O => \N__22731\,
            I => \N__22719\
        );

    \I__2978\ : Span4Mux_h
    port map (
            O => \N__22728\,
            I => \N__22714\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__22725\,
            I => \N__22714\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__22722\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2975\ : Odrv4
    port map (
            O => \N__22719\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__22714\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2973\ : InMux
    port map (
            O => \N__22707\,
            I => \N__22688\
        );

    \I__2972\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22685\
        );

    \I__2971\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22682\
        );

    \I__2970\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22679\
        );

    \I__2969\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22668\
        );

    \I__2968\ : InMux
    port map (
            O => \N__22702\,
            I => \N__22668\
        );

    \I__2967\ : InMux
    port map (
            O => \N__22701\,
            I => \N__22668\
        );

    \I__2966\ : InMux
    port map (
            O => \N__22700\,
            I => \N__22668\
        );

    \I__2965\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22668\
        );

    \I__2964\ : InMux
    port map (
            O => \N__22698\,
            I => \N__22665\
        );

    \I__2963\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22661\
        );

    \I__2962\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22635\
        );

    \I__2961\ : InMux
    port map (
            O => \N__22695\,
            I => \N__22635\
        );

    \I__2960\ : InMux
    port map (
            O => \N__22694\,
            I => \N__22635\
        );

    \I__2959\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22635\
        );

    \I__2958\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22635\
        );

    \I__2957\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22635\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__22688\,
            I => \N__22632\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22621\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__22682\,
            I => \N__22621\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22621\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__22668\,
            I => \N__22621\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__22665\,
            I => \N__22621\
        );

    \I__2950\ : InMux
    port map (
            O => \N__22664\,
            I => \N__22617\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__22661\,
            I => \N__22614\
        );

    \I__2948\ : InMux
    port map (
            O => \N__22660\,
            I => \N__22599\
        );

    \I__2947\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22599\
        );

    \I__2946\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22599\
        );

    \I__2945\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22599\
        );

    \I__2944\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22599\
        );

    \I__2943\ : InMux
    port map (
            O => \N__22655\,
            I => \N__22599\
        );

    \I__2942\ : InMux
    port map (
            O => \N__22654\,
            I => \N__22599\
        );

    \I__2941\ : InMux
    port map (
            O => \N__22653\,
            I => \N__22596\
        );

    \I__2940\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22585\
        );

    \I__2939\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22585\
        );

    \I__2938\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22585\
        );

    \I__2937\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22585\
        );

    \I__2936\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22585\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22582\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__22632\,
            I => \N__22577\
        );

    \I__2933\ : Span4Mux_v
    port map (
            O => \N__22621\,
            I => \N__22577\
        );

    \I__2932\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22574\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22569\
        );

    \I__2930\ : Span4Mux_h
    port map (
            O => \N__22614\,
            I => \N__22569\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__22599\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__22596\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__22585\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__22582\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__22577\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__22574\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__22569\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__2922\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22551\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__22551\,
            I => \N__22548\
        );

    \I__2920\ : Odrv12
    port map (
            O => \N__22548\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__2919\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__22542\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__2917\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22535\
        );

    \I__2916\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22532\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__22535\,
            I => \N__22529\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22524\
        );

    \I__2913\ : Span12Mux_v
    port map (
            O => \N__22529\,
            I => \N__22524\
        );

    \I__2912\ : Odrv12
    port map (
            O => \N__22524\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__2911\ : InMux
    port map (
            O => \N__22521\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__2910\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22515\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__22515\,
            I => \N__22512\
        );

    \I__2908\ : Span4Mux_s1_h
    port map (
            O => \N__22512\,
            I => \N__22508\
        );

    \I__2907\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22505\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__22508\,
            I => \N__22502\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__22505\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2904\ : Odrv4
    port map (
            O => \N__22502\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__2903\ : InMux
    port map (
            O => \N__22497\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__2902\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22491\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__22491\,
            I => \N__22487\
        );

    \I__2900\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22484\
        );

    \I__2899\ : Span4Mux_s1_h
    port map (
            O => \N__22487\,
            I => \N__22481\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22478\
        );

    \I__2897\ : Span4Mux_h
    port map (
            O => \N__22481\,
            I => \N__22475\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__22478\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__22475\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__2894\ : InMux
    port map (
            O => \N__22470\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__2893\ : InMux
    port map (
            O => \N__22467\,
            I => \N__22463\
        );

    \I__2892\ : InMux
    port map (
            O => \N__22466\,
            I => \N__22460\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__22463\,
            I => \N__22457\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22454\
        );

    \I__2889\ : Span4Mux_v
    port map (
            O => \N__22457\,
            I => \N__22451\
        );

    \I__2888\ : Span4Mux_v
    port map (
            O => \N__22454\,
            I => \N__22448\
        );

    \I__2887\ : Sp12to4
    port map (
            O => \N__22451\,
            I => \N__22445\
        );

    \I__2886\ : Span4Mux_h
    port map (
            O => \N__22448\,
            I => \N__22442\
        );

    \I__2885\ : Odrv12
    port map (
            O => \N__22445\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__22442\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__2883\ : InMux
    port map (
            O => \N__22437\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22430\
        );

    \I__2881\ : InMux
    port map (
            O => \N__22433\,
            I => \N__22427\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__22430\,
            I => \N__22424\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__22427\,
            I => \N__22421\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__22424\,
            I => \N__22418\
        );

    \I__2877\ : Span4Mux_v
    port map (
            O => \N__22421\,
            I => \N__22415\
        );

    \I__2876\ : Span4Mux_h
    port map (
            O => \N__22418\,
            I => \N__22412\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__22415\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__22412\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__2873\ : InMux
    port map (
            O => \N__22407\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22400\
        );

    \I__2871\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22397\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__22400\,
            I => \N__22392\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__22397\,
            I => \N__22392\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__22392\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2867\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22385\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22382\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__22385\,
            I => \N__22379\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22376\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__22379\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__22376\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22368\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__22368\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__22365\,
            I => \N__22361\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22356\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22356\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22356\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2855\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22347\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22347\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22347\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2852\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22340\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22337\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22334\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22331\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__22334\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__22331\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2846\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22322\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22319\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22316\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__22319\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__22316\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__22311\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22305\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22305\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\
        );

    \I__2838\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22296\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22301\,
            I => \N__22296\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22293\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__22293\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22290\,
            I => \N__22284\
        );

    \I__2833\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22284\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22284\,
            I => \N__22281\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__22281\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22272\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22272\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__22272\,
            I => \N__22269\
        );

    \I__2827\ : Odrv12
    port map (
            O => \N__22269\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__22266\,
            I => \N__22263\
        );

    \I__2825\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22257\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22257\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__22257\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__22254\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22245\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22245\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__22245\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2818\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22239\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22239\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\
        );

    \I__2816\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22233\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__22233\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__22230\,
            I => \N__22219\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__22229\,
            I => \N__22215\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__22228\,
            I => \N__22211\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__22227\,
            I => \N__22208\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__22226\,
            I => \N__22204\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__22225\,
            I => \N__22200\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__22224\,
            I => \N__22196\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22178\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22178\
        );

    \I__2805\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22178\
        );

    \I__2804\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22178\
        );

    \I__2803\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22178\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22178\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22178\
        );

    \I__2800\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22161\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22161\
        );

    \I__2798\ : InMux
    port map (
            O => \N__22204\,
            I => \N__22161\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22203\,
            I => \N__22161\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22161\
        );

    \I__2795\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22161\
        );

    \I__2794\ : InMux
    port map (
            O => \N__22196\,
            I => \N__22161\
        );

    \I__2793\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22161\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__22194\,
            I => \N__22158\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__22193\,
            I => \N__22154\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__22178\,
            I => \N__22149\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__22161\,
            I => \N__22149\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22158\,
            I => \N__22142\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22142\
        );

    \I__2786\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22142\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__22149\,
            I => \N__22137\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__22142\,
            I => \N__22137\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__22137\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__22134\,
            I => \N__22131\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22125\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__22125\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22118\
        );

    \I__2777\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22114\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22118\,
            I => \N__22111\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22107\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__22114\,
            I => \N__22104\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__22111\,
            I => \N__22101\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22098\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__22107\,
            I => \N__22095\
        );

    \I__2770\ : Span4Mux_v
    port map (
            O => \N__22104\,
            I => \N__22092\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__22101\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__22098\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__22095\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__22092\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22083\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__22080\,
            I => \N__22077\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22073\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22068\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22065\
        );

    \I__2760\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22062\
        );

    \I__2759\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22059\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__22068\,
            I => \N__22056\
        );

    \I__2757\ : Span4Mux_v
    port map (
            O => \N__22065\,
            I => \N__22053\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22050\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__22059\,
            I => \N__22045\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__22056\,
            I => \N__22045\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__22053\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2752\ : Odrv12
    port map (
            O => \N__22050\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__22045\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22038\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22031\
        );

    \I__2748\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22027\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__22031\,
            I => \N__22023\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \N__22020\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__22027\,
            I => \N__22017\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22014\
        );

    \I__2743\ : Span4Mux_v
    port map (
            O => \N__22023\,
            I => \N__22011\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22020\,
            I => \N__22008\
        );

    \I__2741\ : Sp12to4
    port map (
            O => \N__22017\,
            I => \N__22003\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__22003\
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__22011\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22008\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2737\ : Odrv12
    port map (
            O => \N__22003\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2736\ : InMux
    port map (
            O => \N__21996\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__21993\,
            I => \N__21990\
        );

    \I__2734\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21987\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21983\
        );

    \I__2732\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21978\
        );

    \I__2731\ : Span4Mux_v
    port map (
            O => \N__21983\,
            I => \N__21975\
        );

    \I__2730\ : InMux
    port map (
            O => \N__21982\,
            I => \N__21972\
        );

    \I__2729\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21969\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__21978\,
            I => \N__21966\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__21975\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__21972\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__21969\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__21966\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2723\ : InMux
    port map (
            O => \N__21957\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2722\ : InMux
    port map (
            O => \N__21954\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2721\ : InMux
    port map (
            O => \N__21951\,
            I => \N__21948\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21945\
        );

    \I__2719\ : Span4Mux_s3_h
    port map (
            O => \N__21945\,
            I => \N__21942\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__21942\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2717\ : InMux
    port map (
            O => \N__21939\,
            I => \N__21936\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__21936\,
            I => \N__21932\
        );

    \I__2715\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21929\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__21932\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__21929\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2712\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21921\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__21921\,
            I => \N__21917\
        );

    \I__2710\ : InMux
    port map (
            O => \N__21920\,
            I => \N__21914\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__21917\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__21914\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2707\ : InMux
    port map (
            O => \N__21909\,
            I => \N__21906\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__21906\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__2705\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21899\
        );

    \I__2704\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21896\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__21899\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__21896\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__21891\,
            I => \N__21888\
        );

    \I__2700\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21884\
        );

    \I__2699\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21881\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__21884\,
            I => \N__21878\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21875\
        );

    \I__2696\ : Odrv12
    port map (
            O => \N__21878\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__21875\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2694\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__21867\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\
        );

    \I__2692\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21855\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__21860\,
            I => \N__21852\
        );

    \I__2689\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21849\
        );

    \I__2688\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21846\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__21855\,
            I => \N__21843\
        );

    \I__2686\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21840\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__21849\,
            I => \N__21835\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__21846\,
            I => \N__21835\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__21843\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__21840\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__21835\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2680\ : InMux
    port map (
            O => \N__21828\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__21825\,
            I => \N__21821\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__21824\,
            I => \N__21818\
        );

    \I__2677\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21814\
        );

    \I__2676\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21811\
        );

    \I__2675\ : InMux
    port map (
            O => \N__21817\,
            I => \N__21808\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21805\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__21811\,
            I => \N__21799\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__21808\,
            I => \N__21799\
        );

    \I__2671\ : Span4Mux_v
    port map (
            O => \N__21805\,
            I => \N__21796\
        );

    \I__2670\ : InMux
    port map (
            O => \N__21804\,
            I => \N__21793\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__21799\,
            I => \N__21790\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__21796\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__21793\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__21790\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2665\ : InMux
    port map (
            O => \N__21783\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2664\ : InMux
    port map (
            O => \N__21780\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2663\ : InMux
    port map (
            O => \N__21777\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2662\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21770\
        );

    \I__2661\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21765\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__21770\,
            I => \N__21762\
        );

    \I__2659\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21759\
        );

    \I__2658\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21756\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__21765\,
            I => \N__21753\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__21762\,
            I => \N__21750\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__21759\,
            I => \N__21747\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__21756\,
            I => \N__21742\
        );

    \I__2653\ : Span4Mux_v
    port map (
            O => \N__21753\,
            I => \N__21742\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__21750\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2651\ : Odrv12
    port map (
            O => \N__21747\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__21742\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2649\ : InMux
    port map (
            O => \N__21735\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__21732\,
            I => \N__21728\
        );

    \I__2647\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21725\
        );

    \I__2646\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21721\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21717\
        );

    \I__2644\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21714\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__21721\,
            I => \N__21711\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__21720\,
            I => \N__21708\
        );

    \I__2641\ : Span4Mux_h
    port map (
            O => \N__21717\,
            I => \N__21703\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__21714\,
            I => \N__21703\
        );

    \I__2639\ : Span4Mux_v
    port map (
            O => \N__21711\,
            I => \N__21700\
        );

    \I__2638\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21697\
        );

    \I__2637\ : Span4Mux_v
    port map (
            O => \N__21703\,
            I => \N__21694\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__21700\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__21697\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__21694\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__21687\,
            I => \N__21684\
        );

    \I__2632\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21680\
        );

    \I__2631\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21677\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__21680\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__21677\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2628\ : InMux
    port map (
            O => \N__21672\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2627\ : InMux
    port map (
            O => \N__21669\,
            I => \N__21665\
        );

    \I__2626\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21662\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21659\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__21662\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__21659\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2622\ : InMux
    port map (
            O => \N__21654\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__21651\,
            I => \N__21647\
        );

    \I__2620\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21644\
        );

    \I__2619\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21640\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__21644\,
            I => \N__21636\
        );

    \I__2617\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21633\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__21640\,
            I => \N__21630\
        );

    \I__2615\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21627\
        );

    \I__2614\ : Span4Mux_v
    port map (
            O => \N__21636\,
            I => \N__21622\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21622\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__21630\,
            I => \N__21619\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__21627\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__21622\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__21619\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2608\ : InMux
    port map (
            O => \N__21612\,
            I => \bfn_3_20_0_\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__21609\,
            I => \N__21605\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__21608\,
            I => \N__21602\
        );

    \I__2605\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21599\
        );

    \I__2604\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21593\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__21596\,
            I => \N__21588\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__21593\,
            I => \N__21585\
        );

    \I__2600\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21582\
        );

    \I__2599\ : InMux
    port map (
            O => \N__21591\,
            I => \N__21579\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__21588\,
            I => \N__21576\
        );

    \I__2597\ : Sp12to4
    port map (
            O => \N__21585\,
            I => \N__21571\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__21582\,
            I => \N__21571\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__21579\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__21576\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2593\ : Odrv12
    port map (
            O => \N__21571\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2592\ : InMux
    port map (
            O => \N__21564\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2591\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21558\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21555\
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__21555\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__21552\,
            I => \N__21548\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__21551\,
            I => \N__21545\
        );

    \I__2586\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21542\
        );

    \I__2585\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21539\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__21542\,
            I => \N__21536\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__21539\,
            I => \N__21530\
        );

    \I__2582\ : Span4Mux_h
    port map (
            O => \N__21536\,
            I => \N__21530\
        );

    \I__2581\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21526\
        );

    \I__2580\ : Span4Mux_v
    port map (
            O => \N__21530\,
            I => \N__21523\
        );

    \I__2579\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21520\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__21526\,
            I => \N__21517\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__21523\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__21520\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2575\ : Odrv12
    port map (
            O => \N__21517\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2574\ : InMux
    port map (
            O => \N__21510\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2573\ : InMux
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__21501\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__21498\,
            I => \N__21495\
        );

    \I__2569\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21491\
        );

    \I__2568\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21488\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21484\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__21488\,
            I => \N__21481\
        );

    \I__2565\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21478\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__21484\,
            I => \N__21474\
        );

    \I__2563\ : Span12Mux_s2_h
    port map (
            O => \N__21481\,
            I => \N__21469\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__21478\,
            I => \N__21469\
        );

    \I__2561\ : InMux
    port map (
            O => \N__21477\,
            I => \N__21466\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__21474\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2559\ : Odrv12
    port map (
            O => \N__21469\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__21466\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2557\ : InMux
    port map (
            O => \N__21459\,
            I => \N__21455\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21458\,
            I => \N__21452\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__21455\,
            I => \N__21447\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__21452\,
            I => \N__21447\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__21447\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2552\ : InMux
    port map (
            O => \N__21444\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__21441\,
            I => \N__21438\
        );

    \I__2550\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21432\
        );

    \I__2549\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21429\
        );

    \I__2548\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21426\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21423\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__21432\,
            I => \N__21418\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21429\,
            I => \N__21418\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__21426\,
            I => \N__21415\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21412\
        );

    \I__2542\ : Span4Mux_h
    port map (
            O => \N__21418\,
            I => \N__21407\
        );

    \I__2541\ : Span4Mux_h
    port map (
            O => \N__21415\,
            I => \N__21407\
        );

    \I__2540\ : Odrv12
    port map (
            O => \N__21412\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__21407\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2538\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21399\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__21399\,
            I => \N__21395\
        );

    \I__2536\ : InMux
    port map (
            O => \N__21398\,
            I => \N__21392\
        );

    \I__2535\ : Span4Mux_s3_h
    port map (
            O => \N__21395\,
            I => \N__21387\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21387\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__21387\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2532\ : InMux
    port map (
            O => \N__21384\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21378\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__2529\ : Odrv12
    port map (
            O => \N__21375\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__21372\,
            I => \N__21367\
        );

    \I__2527\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21364\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21361\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21357\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21354\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21351\
        );

    \I__2522\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21348\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21357\,
            I => \N__21345\
        );

    \I__2520\ : Span4Mux_s3_h
    port map (
            O => \N__21354\,
            I => \N__21340\
        );

    \I__2519\ : Span4Mux_s3_h
    port map (
            O => \N__21351\,
            I => \N__21340\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21337\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__21345\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__21340\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__21337\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__21330\,
            I => \N__21327\
        );

    \I__2513\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21323\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21320\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__21323\,
            I => \N__21317\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21320\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2509\ : Odrv4
    port map (
            O => \N__21317\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21312\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2507\ : InMux
    port map (
            O => \N__21309\,
            I => \N__21305\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21308\,
            I => \N__21302\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21297\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__21302\,
            I => \N__21294\
        );

    \I__2503\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21291\
        );

    \I__2502\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21288\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__21297\,
            I => \N__21283\
        );

    \I__2500\ : Span4Mux_h
    port map (
            O => \N__21294\,
            I => \N__21283\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21291\,
            I => \N__21278\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__21288\,
            I => \N__21278\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__21283\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__21278\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2495\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21269\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21272\,
            I => \N__21266\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__21269\,
            I => \N__21263\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__21266\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__21263\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2490\ : InMux
    port map (
            O => \N__21258\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__21255\,
            I => \N__21252\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21248\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21244\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__21248\,
            I => \N__21240\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21237\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21234\
        );

    \I__2483\ : InMux
    port map (
            O => \N__21243\,
            I => \N__21231\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__21240\,
            I => \N__21228\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__21237\,
            I => \N__21225\
        );

    \I__2480\ : Sp12to4
    port map (
            O => \N__21234\,
            I => \N__21220\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21220\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__21228\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__21225\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2476\ : Odrv12
    port map (
            O => \N__21220\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2475\ : InMux
    port map (
            O => \N__21213\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__21210\,
            I => \N__21205\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21202\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21199\
        );

    \I__2471\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21196\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21192\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21189\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21186\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21183\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__21192\,
            I => \N__21180\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21175\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__21186\,
            I => \N__21175\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21183\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__21180\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__21175\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21168\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__2458\ : InMux
    port map (
            O => \N__21162\,
            I => \N__21157\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__21161\,
            I => \N__21154\
        );

    \I__2456\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21151\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__21157\,
            I => \N__21148\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21145\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21151\,
            I => \N__21142\
        );

    \I__2452\ : Span4Mux_h
    port map (
            O => \N__21148\,
            I => \N__21136\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__21145\,
            I => \N__21136\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__21142\,
            I => \N__21133\
        );

    \I__2449\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21130\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__21136\,
            I => \N__21127\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__21133\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21130\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__21127\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21120\,
            I => \bfn_3_19_0_\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__21111\
        );

    \I__2441\ : Odrv12
    port map (
            O => \N__21111\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__21108\,
            I => \N__21103\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21098\
        );

    \I__2438\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21098\
        );

    \I__2437\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21095\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__21098\,
            I => \N__21091\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21088\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__21094\,
            I => \N__21085\
        );

    \I__2433\ : Span4Mux_v
    port map (
            O => \N__21091\,
            I => \N__21082\
        );

    \I__2432\ : Span4Mux_v
    port map (
            O => \N__21088\,
            I => \N__21079\
        );

    \I__2431\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21076\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__21082\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__21079\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__21076\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2427\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21066\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21061\
        );

    \I__2425\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21056\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21056\
        );

    \I__2423\ : Span4Mux_v
    port map (
            O => \N__21061\,
            I => \N__21051\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__21051\
        );

    \I__2421\ : Span4Mux_v
    port map (
            O => \N__21051\,
            I => \N__21048\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__21048\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21045\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2418\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21039\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21039\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__21036\,
            I => \N__21031\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21026\
        );

    \I__2414\ : InMux
    port map (
            O => \N__21034\,
            I => \N__21026\
        );

    \I__2413\ : InMux
    port map (
            O => \N__21031\,
            I => \N__21023\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__21026\,
            I => \N__21017\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__21023\,
            I => \N__21017\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21014\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__21017\,
            I => \N__21011\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__21008\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__21011\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__21008\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2405\ : InMux
    port map (
            O => \N__21003\,
            I => \N__20999\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20996\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20989\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__20996\,
            I => \N__20989\
        );

    \I__2401\ : InMux
    port map (
            O => \N__20995\,
            I => \N__20984\
        );

    \I__2400\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20984\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__20989\,
            I => \N__20979\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__20984\,
            I => \N__20979\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__20979\,
            I => \N__20976\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__20976\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2395\ : InMux
    port map (
            O => \N__20973\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2394\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20967\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__20967\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__20964\,
            I => \N__20961\
        );

    \I__2391\ : InMux
    port map (
            O => \N__20961\,
            I => \N__20958\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__20958\,
            I => \N__20953\
        );

    \I__2389\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20948\
        );

    \I__2388\ : InMux
    port map (
            O => \N__20956\,
            I => \N__20948\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__20953\,
            I => \N__20943\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__20948\,
            I => \N__20943\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__20943\,
            I => \N__20939\
        );

    \I__2384\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20936\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__20939\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__20936\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2381\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20928\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__20928\,
            I => \N__20923\
        );

    \I__2379\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20920\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__20926\,
            I => \N__20917\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__20923\,
            I => \N__20914\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20911\
        );

    \I__2375\ : InMux
    port map (
            O => \N__20917\,
            I => \N__20908\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__20914\,
            I => \N__20905\
        );

    \I__2373\ : Span4Mux_v
    port map (
            O => \N__20911\,
            I => \N__20900\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__20908\,
            I => \N__20900\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__20905\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__20900\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2369\ : InMux
    port map (
            O => \N__20895\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2368\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20886\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__20886\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__20883\,
            I => \N__20879\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__20882\,
            I => \N__20875\
        );

    \I__2363\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20872\
        );

    \I__2362\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20869\
        );

    \I__2361\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20866\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__20872\,
            I => \N__20863\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20857\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20857\
        );

    \I__2357\ : Span4Mux_v
    port map (
            O => \N__20863\,
            I => \N__20854\
        );

    \I__2356\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20851\
        );

    \I__2355\ : Odrv12
    port map (
            O => \N__20857\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__20854\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__20851\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2352\ : InMux
    port map (
            O => \N__20844\,
            I => \N__20841\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__20841\,
            I => \N__20837\
        );

    \I__2350\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20834\
        );

    \I__2349\ : Span4Mux_s3_h
    port map (
            O => \N__20837\,
            I => \N__20830\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__20834\,
            I => \N__20827\
        );

    \I__2347\ : InMux
    port map (
            O => \N__20833\,
            I => \N__20824\
        );

    \I__2346\ : Span4Mux_v
    port map (
            O => \N__20830\,
            I => \N__20821\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__20827\,
            I => \N__20816\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__20824\,
            I => \N__20816\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__20821\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__20816\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2341\ : InMux
    port map (
            O => \N__20811\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2340\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__20805\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \N__20799\
        );

    \I__2337\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20792\
        );

    \I__2335\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20787\
        );

    \I__2334\ : Span4Mux_h
    port map (
            O => \N__20792\,
            I => \N__20784\
        );

    \I__2333\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20779\
        );

    \I__2332\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20779\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__20787\,
            I => \N__20776\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__20784\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__20779\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2328\ : Odrv12
    port map (
            O => \N__20776\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__2326\ : InMux
    port map (
            O => \N__20766\,
            I => \N__20761\
        );

    \I__2325\ : InMux
    port map (
            O => \N__20765\,
            I => \N__20758\
        );

    \I__2324\ : InMux
    port map (
            O => \N__20764\,
            I => \N__20755\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__20761\,
            I => \N__20752\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20749\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__20755\,
            I => \N__20746\
        );

    \I__2320\ : Span12Mux_s3_h
    port map (
            O => \N__20752\,
            I => \N__20743\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__20749\,
            I => \N__20738\
        );

    \I__2318\ : Span4Mux_s3_h
    port map (
            O => \N__20746\,
            I => \N__20738\
        );

    \I__2317\ : Odrv12
    port map (
            O => \N__20743\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__20738\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2315\ : InMux
    port map (
            O => \N__20733\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__20730\,
            I => \N__20724\
        );

    \I__2313\ : InMux
    port map (
            O => \N__20729\,
            I => \N__20719\
        );

    \I__2312\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20719\
        );

    \I__2311\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20716\
        );

    \I__2310\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20713\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__20719\,
            I => \N__20710\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20707\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20704\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__20710\,
            I => \N__20701\
        );

    \I__2305\ : Span4Mux_s3_h
    port map (
            O => \N__20707\,
            I => \N__20698\
        );

    \I__2304\ : Odrv12
    port map (
            O => \N__20704\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__20701\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__20698\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2301\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20684\
        );

    \I__2299\ : InMux
    port map (
            O => \N__20687\,
            I => \N__20680\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__20684\,
            I => \N__20677\
        );

    \I__2297\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20674\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20671\
        );

    \I__2295\ : Span4Mux_v
    port map (
            O => \N__20677\,
            I => \N__20668\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__20674\,
            I => \N__20663\
        );

    \I__2293\ : Span4Mux_v
    port map (
            O => \N__20671\,
            I => \N__20663\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__20668\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__20663\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2290\ : InMux
    port map (
            O => \N__20658\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__2289\ : CascadeMux
    port map (
            O => \N__20655\,
            I => \N__20651\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \N__20648\
        );

    \I__2287\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20643\
        );

    \I__2286\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20640\
        );

    \I__2285\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20635\
        );

    \I__2284\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20635\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__20643\,
            I => \N__20632\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__20640\,
            I => \N__20629\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__20635\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__20632\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__20629\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__20622\,
            I => \N__20619\
        );

    \I__2277\ : InMux
    port map (
            O => \N__20619\,
            I => \N__20616\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20612\
        );

    \I__2275\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20609\
        );

    \I__2274\ : Span4Mux_s3_h
    port map (
            O => \N__20612\,
            I => \N__20605\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20602\
        );

    \I__2272\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20599\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__20605\,
            I => \N__20596\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__20602\,
            I => \N__20591\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__20599\,
            I => \N__20591\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__20596\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__20591\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2266\ : InMux
    port map (
            O => \N__20586\,
            I => \bfn_3_18_0_\
        );

    \I__2265\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20580\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__20580\,
            I => \N__20577\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__20577\,
            I => \N__20574\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__20574\,
            I => \N__20571\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__20571\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__2260\ : InMux
    port map (
            O => \N__20568\,
            I => \N__20562\
        );

    \I__2259\ : InMux
    port map (
            O => \N__20567\,
            I => \N__20548\
        );

    \I__2258\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20545\
        );

    \I__2257\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20542\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20539\
        );

    \I__2255\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20536\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__20560\,
            I => \N__20533\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__20559\,
            I => \N__20530\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__20558\,
            I => \N__20527\
        );

    \I__2251\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20508\
        );

    \I__2250\ : InMux
    port map (
            O => \N__20556\,
            I => \N__20505\
        );

    \I__2249\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20494\
        );

    \I__2248\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20494\
        );

    \I__2247\ : InMux
    port map (
            O => \N__20553\,
            I => \N__20494\
        );

    \I__2246\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20494\
        );

    \I__2245\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20494\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__20548\,
            I => \N__20483\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__20545\,
            I => \N__20483\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20483\
        );

    \I__2241\ : Span4Mux_h
    port map (
            O => \N__20539\,
            I => \N__20483\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__20536\,
            I => \N__20483\
        );

    \I__2239\ : InMux
    port map (
            O => \N__20533\,
            I => \N__20470\
        );

    \I__2238\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20470\
        );

    \I__2237\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20470\
        );

    \I__2236\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20470\
        );

    \I__2235\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20470\
        );

    \I__2234\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20470\
        );

    \I__2233\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20467\
        );

    \I__2232\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20452\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20452\
        );

    \I__2230\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20452\
        );

    \I__2229\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20452\
        );

    \I__2228\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20452\
        );

    \I__2227\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20452\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20452\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20441\
        );

    \I__2224\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20441\
        );

    \I__2223\ : InMux
    port map (
            O => \N__20513\,
            I => \N__20441\
        );

    \I__2222\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20441\
        );

    \I__2221\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20441\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20434\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20434\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__20494\,
            I => \N__20434\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__20483\,
            I => \N__20431\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20422\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20422\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__20452\,
            I => \N__20422\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__20441\,
            I => \N__20422\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__20434\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__20431\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__20422\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__20415\,
            I => \N__20412\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20409\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__20409\,
            I => \N__20406\
        );

    \I__2206\ : Span4Mux_h
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__20403\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__20400\,
            I => \N__20391\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__20399\,
            I => \N__20388\
        );

    \I__2202\ : InMux
    port map (
            O => \N__20398\,
            I => \N__20382\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20397\,
            I => \N__20379\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20357\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20357\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20357\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20391\,
            I => \N__20357\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20357\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20387\,
            I => \N__20347\
        );

    \I__2194\ : InMux
    port map (
            O => \N__20386\,
            I => \N__20344\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20341\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__20382\,
            I => \N__20336\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__20379\,
            I => \N__20336\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20333\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20326\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20326\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20326\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20317\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20317\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20317\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20317\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__20370\,
            I => \N__20311\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__20369\,
            I => \N__20308\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__20368\,
            I => \N__20305\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__20357\,
            I => \N__20302\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20287\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20287\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20287\
        );

    \I__2175\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20287\
        );

    \I__2174\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20287\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20287\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20287\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__20347\,
            I => \N__20282\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__20344\,
            I => \N__20282\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__20341\,
            I => \N__20277\
        );

    \I__2168\ : Span4Mux_v
    port map (
            O => \N__20336\,
            I => \N__20277\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20333\,
            I => \N__20274\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20269\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20269\
        );

    \I__2164\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20266\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20315\,
            I => \N__20255\
        );

    \I__2162\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20255\
        );

    \I__2161\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20255\
        );

    \I__2160\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20255\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20255\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__20302\,
            I => \N__20250\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20250\
        );

    \I__2156\ : Span4Mux_v
    port map (
            O => \N__20282\,
            I => \N__20245\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__20277\,
            I => \N__20245\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__20274\,
            I => \N__20240\
        );

    \I__2153\ : Span4Mux_v
    port map (
            O => \N__20269\,
            I => \N__20240\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20266\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20255\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__20250\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__20245\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__20240\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20225\
        );

    \I__2146\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20222\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20219\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__20222\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__20219\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__20214\,
            I => \N__20210\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20206\
        );

    \I__2140\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20203\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__20209\,
            I => \N__20200\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__20206\,
            I => \N__20195\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__20203\,
            I => \N__20195\
        );

    \I__2136\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20191\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__20195\,
            I => \N__20188\
        );

    \I__2134\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20184\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__20191\,
            I => \N__20181\
        );

    \I__2132\ : Span4Mux_s3_h
    port map (
            O => \N__20188\,
            I => \N__20178\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20187\,
            I => \N__20175\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20184\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__20181\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__20178\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__20175\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__20166\,
            I => \N__20162\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20159\
        );

    \I__2124\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20156\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__20159\,
            I => \N__20152\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20156\,
            I => \N__20149\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20146\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__20152\,
            I => \N__20143\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__20149\,
            I => \N__20140\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20146\,
            I => \N__20137\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__20143\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2116\ : Odrv4
    port map (
            O => \N__20140\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__20137\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20127\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20127\,
            I => \N__20124\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__20121\,
            I => \N__20118\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__20118\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20115\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2108\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20109\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__20109\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\
        );

    \I__2106\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20102\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20098\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20102\,
            I => \N__20095\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20092\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20098\,
            I => \N__20089\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__20095\,
            I => pwm_duty_input_4
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20092\,
            I => pwm_duty_input_4
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__20089\,
            I => pwm_duty_input_4
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__20082\,
            I => \N__20079\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20075\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20071\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20075\,
            I => \N__20068\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20065\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20071\,
            I => \N__20062\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__20068\,
            I => pwm_duty_input_3
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__20065\,
            I => pwm_duty_input_3
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__20062\,
            I => pwm_duty_input_3
        );

    \I__2089\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20051\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20048\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__20044\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20048\,
            I => \N__20041\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20038\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__20044\,
            I => \N__20035\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__20041\,
            I => pwm_duty_input_5
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__20038\,
            I => pwm_duty_input_5
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__20035\,
            I => pwm_duty_input_5
        );

    \I__2080\ : InMux
    port map (
            O => \N__20028\,
            I => \N__20025\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__20022\,
            I => \rgb_drv_RNOZ0\
        );

    \I__2077\ : InMux
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__20016\,
            I => \N__20013\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__20013\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__20010\,
            I => \N__20007\
        );

    \I__2073\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__20001\,
            I => \N__19998\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__19998\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__2068\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19989\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__19989\,
            I => \N__19986\
        );

    \I__2066\ : Span4Mux_h
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__19983\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__19980\,
            I => \N__19977\
        );

    \I__2063\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19971\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__19971\,
            I => \N__19968\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__19968\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__19965\,
            I => \N__19957\
        );

    \I__2058\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19948\
        );

    \I__2057\ : InMux
    port map (
            O => \N__19963\,
            I => \N__19948\
        );

    \I__2056\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19948\
        );

    \I__2055\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19948\
        );

    \I__2054\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19940\
        );

    \I__2053\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19940\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19937\
        );

    \I__2051\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19934\
        );

    \I__2050\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19931\
        );

    \I__2049\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19928\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__19940\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__19937\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__19934\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__19931\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__19928\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__19917\,
            I => \N__19914\
        );

    \I__2042\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19908\
        );

    \I__2041\ : InMux
    port map (
            O => \N__19913\,
            I => \N__19908\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__19908\,
            I => \N__19904\
        );

    \I__2039\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19901\
        );

    \I__2038\ : Odrv12
    port map (
            O => \N__19904\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__19901\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2036\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__19893\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__19890\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\
        );

    \I__2033\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19883\
        );

    \I__2032\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19880\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__19883\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__19880\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2029\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19872\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19868\
        );

    \I__2027\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19865\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__19868\,
            I => \N__19862\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__19865\,
            I => pwm_duty_input_0
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__19862\,
            I => pwm_duty_input_0
        );

    \I__2023\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19853\
        );

    \I__2022\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19850\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__19853\,
            I => \N__19847\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__19850\,
            I => pwm_duty_input_1
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__19847\,
            I => pwm_duty_input_1
        );

    \I__2018\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__19839\,
            I => \N__19835\
        );

    \I__2016\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19832\
        );

    \I__2015\ : Span4Mux_s1_h
    port map (
            O => \N__19835\,
            I => \N__19829\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__19832\,
            I => pwm_duty_input_2
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__19829\,
            I => pwm_duty_input_2
        );

    \I__2012\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19819\
        );

    \I__2011\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19814\
        );

    \I__2010\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19814\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__19819\,
            I => \N__19811\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__19814\,
            I => pwm_duty_input_7
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__19811\,
            I => pwm_duty_input_7
        );

    \I__2006\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19803\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19798\
        );

    \I__2004\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19793\
        );

    \I__2003\ : InMux
    port map (
            O => \N__19801\,
            I => \N__19793\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__19798\,
            I => \N__19790\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__19793\,
            I => pwm_duty_input_8
        );

    \I__2000\ : Odrv4
    port map (
            O => \N__19790\,
            I => pwm_duty_input_8
        );

    \I__1999\ : InMux
    port map (
            O => \N__19785\,
            I => \N__19781\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__19784\,
            I => \N__19777\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__19781\,
            I => \N__19774\
        );

    \I__1996\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19769\
        );

    \I__1995\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19769\
        );

    \I__1994\ : Span4Mux_s1_h
    port map (
            O => \N__19774\,
            I => \N__19766\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__19769\,
            I => pwm_duty_input_6
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__19766\,
            I => pwm_duty_input_6
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__19761\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\
        );

    \I__1990\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__19755\,
            I => \N__19750\
        );

    \I__1988\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19745\
        );

    \I__1987\ : InMux
    port map (
            O => \N__19753\,
            I => \N__19745\
        );

    \I__1986\ : Span4Mux_s1_h
    port map (
            O => \N__19750\,
            I => \N__19742\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__19745\,
            I => pwm_duty_input_9
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__19742\,
            I => pwm_duty_input_9
        );

    \I__1983\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__19734\,
            I => \pwm_generator_inst.un1_duty_inputlt3\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__19731\,
            I => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__19728\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\
        );

    \I__1979\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__19722\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\
        );

    \I__1977\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__19716\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__19713\,
            I => \N__19710\
        );

    \I__1974\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19707\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__19707\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__19704\,
            I => \N__19696\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__19703\,
            I => \N__19693\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__19702\,
            I => \N__19690\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__19701\,
            I => \N__19687\
        );

    \I__1968\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19678\
        );

    \I__1967\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19678\
        );

    \I__1966\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19678\
        );

    \I__1965\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19678\
        );

    \I__1964\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19674\
        );

    \I__1963\ : InMux
    port map (
            O => \N__19687\,
            I => \N__19671\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__19678\,
            I => \N__19668\
        );

    \I__1961\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19665\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__19674\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__19671\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__19668\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__19665\,
            I => \current_shift_inst.PI_CTRL.N_159\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__19656\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\
        );

    \I__1955\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19650\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__19650\,
            I => \N__19647\
        );

    \I__1953\ : Odrv4
    port map (
            O => \N__19647\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__19644\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\
        );

    \I__1951\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19632\
        );

    \I__1950\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19632\
        );

    \I__1949\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19632\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__19632\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__19629\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__19626\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\
        );

    \I__1945\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__19620\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__1943\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19614\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__19614\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__19611\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\
        );

    \I__1940\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19605\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__19605\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__1938\ : InMux
    port map (
            O => \N__19602\,
            I => \N__19599\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__19599\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__19596\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1935\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__19590\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__1932\ : InMux
    port map (
            O => \N__19584\,
            I => \N__19581\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__19581\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__1930\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__19575\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__19572\,
            I => \N__19569\
        );

    \I__1927\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__19560\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__19557\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__19554\,
            I => \current_shift_inst.PI_CTRL.N_77_cascade_\
        );

    \I__1921\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__19548\,
            I => \current_shift_inst.PI_CTRL.N_43\
        );

    \I__1919\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19542\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__19542\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\
        );

    \I__1917\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__19536\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1914\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19527\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__19527\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__1912\ : InMux
    port map (
            O => \N__19524\,
            I => \N__19521\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__19521\,
            I => \N__19518\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__19518\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__1908\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__19509\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__19506\,
            I => \N__19503\
        );

    \I__1905\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19500\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__19500\,
            I => \N__19497\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__19497\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__19494\,
            I => \N__19491\
        );

    \I__1901\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19488\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__19488\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__1898\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19479\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__19479\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__19476\,
            I => \N__19473\
        );

    \I__1895\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__19470\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__1893\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__19464\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__1891\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N_38_i_i\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__19455\,
            I => \N__19451\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__19454\,
            I => \N__19448\
        );

    \I__1887\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19445\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19442\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__19445\,
            I => \N__19437\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19437\
        );

    \I__1883\ : Span4Mux_v
    port map (
            O => \N__19437\,
            I => \N__19434\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__19434\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__19431\,
            I => \N__19428\
        );

    \I__1880\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19425\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__19425\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19419\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19419\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19413\,
            I => \N__19410\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19410\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__1872\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19401\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__19398\,
            I => \N__19395\
        );

    \I__1869\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__19392\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__19389\,
            I => \N__19386\
        );

    \I__1866\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19383\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__19383\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__19380\,
            I => \N__19377\
        );

    \I__1863\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19374\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__19374\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__19371\,
            I => \N__19367\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__19370\,
            I => \N__19364\
        );

    \I__1859\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19358\
        );

    \I__1858\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19358\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__19363\,
            I => \N__19355\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__19358\,
            I => \N__19352\
        );

    \I__1855\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19349\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__19352\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__19349\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_3\
        );

    \I__1852\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19340\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19337\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__19340\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__19337\,
            I => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19320\
        );

    \I__1847\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19320\
        );

    \I__1846\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19320\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19320\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__19320\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__19317\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19311\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__19311\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__19308\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__19302\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19296\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19296\,
            I => \N__19293\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__19293\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__19290\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__19287\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__19281\,
            I => \N__19278\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__19278\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__19275\,
            I => \N__19272\
        );

    \I__1828\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19269\,
            I => \N__19266\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__19266\,
            I => \N__19263\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__19263\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__1824\ : InMux
    port map (
            O => \N__19260\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__1823\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19254\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__19254\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__1821\ : InMux
    port map (
            O => \N__19251\,
            I => \N__19248\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__19248\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__19245\,
            I => \N__19242\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19239\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19239\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__1816\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__1814\ : Odrv12
    port map (
            O => \N__19230\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19221\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19218\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__19218\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\
        );

    \I__1808\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19209\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__19209\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19200\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__19200\,
            I => \N__19197\
        );

    \I__1803\ : Odrv12
    port map (
            O => \N__19197\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1802\ : InMux
    port map (
            O => \N__19194\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19188\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__19188\,
            I => \N__19185\
        );

    \I__1799\ : Odrv12
    port map (
            O => \N__19185\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19182\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__19179\,
            I => \N__19176\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19173\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__19173\,
            I => \N__19170\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__19170\,
            I => \N__19167\
        );

    \I__1793\ : Odrv4
    port map (
            O => \N__19167\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19164\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__19161\,
            I => \N__19158\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19155\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19152\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__19149\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__1786\ : InMux
    port map (
            O => \N__19146\,
            I => \bfn_1_15_0_\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__1784\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19137\,
            I => \N__19134\
        );

    \I__1782\ : Odrv12
    port map (
            O => \N__19134\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__1781\ : InMux
    port map (
            O => \N__19131\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__19128\,
            I => \N__19125\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19122\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__19122\,
            I => \N__19119\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__19119\,
            I => \N__19116\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__19116\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__1775\ : InMux
    port map (
            O => \N__19113\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__19110\,
            I => \N__19107\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19104\,
            I => \N__19101\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__19101\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19098\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19092\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__19092\,
            I => \N__19089\
        );

    \I__1767\ : Odrv12
    port map (
            O => \N__19089\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19086\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__19083\,
            I => \N__19080\
        );

    \I__1764\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19077\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__19077\,
            I => \N__19074\
        );

    \I__1762\ : Span4Mux_v
    port map (
            O => \N__19074\,
            I => \N__19071\
        );

    \I__1761\ : Odrv4
    port map (
            O => \N__19071\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19068\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__19065\,
            I => \N__19062\
        );

    \I__1758\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19059\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19059\,
            I => \N__19056\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__19056\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19053\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__19050\,
            I => \N__19047\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19044\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19041\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__19041\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1750\ : InMux
    port map (
            O => \N__19038\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__19035\,
            I => \N__19032\
        );

    \I__1748\ : InMux
    port map (
            O => \N__19032\,
            I => \N__19029\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__19029\,
            I => \N__19026\
        );

    \I__1746\ : Span4Mux_v
    port map (
            O => \N__19026\,
            I => \N__19023\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__19023\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19020\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19014\,
            I => \N__19011\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19011\,
            I => \N__19008\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__19005\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19002\,
            I => \bfn_1_14_0_\
        );

    \I__1737\ : InMux
    port map (
            O => \N__18999\,
            I => \N__18996\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__18996\,
            I => \N__18993\
        );

    \I__1735\ : Odrv12
    port map (
            O => \N__18993\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1734\ : InMux
    port map (
            O => \N__18990\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__1732\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18981\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__18981\,
            I => \N__18978\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__18978\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1729\ : InMux
    port map (
            O => \N__18975\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__18972\,
            I => \N__18969\
        );

    \I__1727\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18966\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__18966\,
            I => \N__18963\
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__18963\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1724\ : InMux
    port map (
            O => \N__18960\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__18957\,
            I => \N__18954\
        );

    \I__1722\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__18951\,
            I => \N__18948\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__18948\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1719\ : InMux
    port map (
            O => \N__18945\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1718\ : InMux
    port map (
            O => \N__18942\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__18939\,
            I => \N__18936\
        );

    \I__1716\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18933\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__18930\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1713\ : InMux
    port map (
            O => \N__18927\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__18924\,
            I => \N__18921\
        );

    \I__1711\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18918\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__18918\,
            I => \N__18915\
        );

    \I__1709\ : Span4Mux_h
    port map (
            O => \N__18915\,
            I => \N__18912\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__18912\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1707\ : InMux
    port map (
            O => \N__18909\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__1705\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18900\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__18900\,
            I => \N__18897\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__18897\,
            I => \N__18894\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__18894\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1701\ : InMux
    port map (
            O => \N__18891\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1700\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18885\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__18882\,
            I => \N__18879\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__18879\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1696\ : InMux
    port map (
            O => \N__18876\,
            I => \bfn_1_13_0_\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \N__18870\
        );

    \I__1694\ : InMux
    port map (
            O => \N__18870\,
            I => \N__18867\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__18867\,
            I => \N__18864\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__18864\,
            I => \N__18861\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__18861\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1690\ : InMux
    port map (
            O => \N__18858\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__18855\,
            I => \N__18852\
        );

    \I__1688\ : InMux
    port map (
            O => \N__18852\,
            I => \N__18849\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__18849\,
            I => \N__18846\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__18846\,
            I => \N__18843\
        );

    \I__1685\ : Span4Mux_s1_h
    port map (
            O => \N__18843\,
            I => \N__18840\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__18840\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1683\ : InMux
    port map (
            O => \N__18837\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__18834\,
            I => \N__18831\
        );

    \I__1681\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18828\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__18828\,
            I => \N__18825\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__18825\,
            I => \N__18822\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__18822\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1677\ : InMux
    port map (
            O => \N__18819\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__18816\,
            I => \N__18813\
        );

    \I__1675\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18810\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__18810\,
            I => \N__18807\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__18807\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1672\ : InMux
    port map (
            O => \N__18804\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1671\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18798\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__18798\,
            I => \N__18795\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__18795\,
            I => \N__18792\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__18792\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1667\ : InMux
    port map (
            O => \N__18789\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1666\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__18783\,
            I => \N__18780\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__18780\,
            I => \N__18777\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__18777\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1662\ : InMux
    port map (
            O => \N__18774\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1661\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18768\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__18765\,
            I => \N__18762\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__18762\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__18759\,
            I => \N__18754\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__18758\,
            I => \N__18750\
        );

    \I__1655\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18741\
        );

    \I__1654\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18741\
        );

    \I__1653\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18741\
        );

    \I__1652\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18741\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__18741\,
            I => \N__18730\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__18740\,
            I => \N__18727\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__18739\,
            I => \N__18724\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__18738\,
            I => \N__18721\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__18737\,
            I => \N__18718\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__18736\,
            I => \N__18715\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__18735\,
            I => \N__18712\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__18734\,
            I => \N__18709\
        );

    \I__1643\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18706\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__18730\,
            I => \N__18703\
        );

    \I__1641\ : InMux
    port map (
            O => \N__18727\,
            I => \N__18696\
        );

    \I__1640\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18696\
        );

    \I__1639\ : InMux
    port map (
            O => \N__18721\,
            I => \N__18696\
        );

    \I__1638\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18687\
        );

    \I__1637\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18687\
        );

    \I__1636\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18687\
        );

    \I__1635\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18687\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18682\
        );

    \I__1633\ : Span4Mux_s1_h
    port map (
            O => \N__18703\,
            I => \N__18682\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__18696\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__18687\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__18682\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1629\ : InMux
    port map (
            O => \N__18675\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1628\ : InMux
    port map (
            O => \N__18672\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__18669\,
            I => \N__18666\
        );

    \I__1626\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__18663\,
            I => \N__18660\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__18660\,
            I => \N__18657\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__18657\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1622\ : InMux
    port map (
            O => \N__18654\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1621\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18648\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__18648\,
            I => \N__18645\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__18645\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1618\ : InMux
    port map (
            O => \N__18642\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__18639\,
            I => \N__18636\
        );

    \I__1616\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18633\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__18633\,
            I => \N__18630\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__18630\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1613\ : InMux
    port map (
            O => \N__18627\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__18624\,
            I => \N__18621\
        );

    \I__1611\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18618\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__18618\,
            I => \N__18615\
        );

    \I__1609\ : Span4Mux_h
    port map (
            O => \N__18615\,
            I => \N__18612\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__18612\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1607\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18606\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18603\
        );

    \I__1605\ : Span4Mux_v
    port map (
            O => \N__18603\,
            I => \N__18600\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__18600\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1603\ : InMux
    port map (
            O => \N__18597\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__18594\,
            I => \N__18591\
        );

    \I__1601\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18588\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__18588\,
            I => \N__18585\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__18582\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1597\ : InMux
    port map (
            O => \N__18579\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1596\ : InMux
    port map (
            O => \N__18576\,
            I => \N__18573\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__18573\,
            I => \N__18570\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__18570\,
            I => \N__18567\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__18567\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1592\ : InMux
    port map (
            O => \N__18564\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__1590\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18555\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__18555\,
            I => \N__18552\
        );

    \I__1588\ : Span4Mux_v
    port map (
            O => \N__18552\,
            I => \N__18549\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__18549\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1586\ : InMux
    port map (
            O => \N__18546\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1585\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18540\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__18540\,
            I => \N__18537\
        );

    \I__1583\ : Span4Mux_v
    port map (
            O => \N__18537\,
            I => \N__18534\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__18534\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1581\ : InMux
    port map (
            O => \N__18531\,
            I => \bfn_1_11_0_\
        );

    \I__1580\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18525\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__18525\,
            I => \N__18522\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__18522\,
            I => \N__18519\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__18519\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1576\ : InMux
    port map (
            O => \N__18516\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1575\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18510\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__18510\,
            I => \N__18507\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__18507\,
            I => \N__18504\
        );

    \I__1572\ : Span4Mux_s1_h
    port map (
            O => \N__18504\,
            I => \N__18501\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__18501\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1570\ : InMux
    port map (
            O => \N__18498\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1569\ : InMux
    port map (
            O => \N__18495\,
            I => \N__18492\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__18492\,
            I => \N__18489\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__18489\,
            I => \N__18486\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__18486\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1565\ : InMux
    port map (
            O => \N__18483\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1564\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18477\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__18477\,
            I => \N__18474\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__18474\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1561\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18468\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__18468\,
            I => \N__18465\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__18465\,
            I => \N__18462\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__18462\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \N__18456\
        );

    \I__1556\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18453\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__18453\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1554\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18447\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__18447\,
            I => \N__18444\
        );

    \I__1552\ : Span4Mux_v
    port map (
            O => \N__18444\,
            I => \N__18441\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__18441\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__18438\,
            I => \N__18435\
        );

    \I__1549\ : InMux
    port map (
            O => \N__18435\,
            I => \N__18432\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__18432\,
            I => \N__18429\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__18429\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1546\ : InMux
    port map (
            O => \N__18426\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1545\ : InMux
    port map (
            O => \N__18423\,
            I => \N__18420\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__18420\,
            I => \N__18417\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__18417\,
            I => \N__18414\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__18414\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__18411\,
            I => \N__18408\
        );

    \I__1540\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18405\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__18405\,
            I => \N__18402\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__18402\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1537\ : InMux
    port map (
            O => \N__18399\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1536\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18393\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__18393\,
            I => \N__18390\
        );

    \I__1534\ : Span4Mux_v
    port map (
            O => \N__18390\,
            I => \N__18387\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__18387\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__1531\ : InMux
    port map (
            O => \N__18381\,
            I => \N__18378\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__18375\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1528\ : InMux
    port map (
            O => \N__18372\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1527\ : IoInMux
    port map (
            O => \N__18369\,
            I => \N__18366\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__1525\ : Span4Mux_s3_v
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__1524\ : Span4Mux_h
    port map (
            O => \N__18360\,
            I => \N__18357\
        );

    \I__1523\ : Sp12to4
    port map (
            O => \N__18357\,
            I => \N__18354\
        );

    \I__1522\ : Span12Mux_s9_v
    port map (
            O => \N__18354\,
            I => \N__18351\
        );

    \I__1521\ : Span12Mux_v
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__1520\ : Odrv12
    port map (
            O => \N__18348\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1519\ : IoInMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18339\
        );

    \I__1517\ : IoSpan4Mux
    port map (
            O => \N__18339\,
            I => \N__18336\
        );

    \I__1516\ : IoSpan4Mux
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__18333\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_16_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_16_14_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_12_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_12_18_0_\
        );

    \IN_MUX_bfv_12_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_12_19_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_14_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_14_20_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_10_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_26_0_\
        );

    \IN_MUX_bfv_10_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_10_27_0_\
        );

    \IN_MUX_bfv_10_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_10_28_0_\
        );

    \IN_MUX_bfv_11_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_24_0_\
        );

    \IN_MUX_bfv_11_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_11_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_7_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_7_28_0_\
        );

    \IN_MUX_bfv_13_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_24_0_\
        );

    \IN_MUX_bfv_13_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_13_25_0_\
        );

    \IN_MUX_bfv_13_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_22_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_13_23_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_12_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_7_0_\
        );

    \IN_MUX_bfv_12_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_12_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_15_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_15_15_0_\
        );

    \IN_MUX_bfv_15_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_15_16_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_17_20_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_5_16_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18369\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18345\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33000\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_162_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__42123\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32487\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__35640\,
            CLKHFEN => \N__35642\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__35641\,
            RGB2PWM => \N__19461\,
            RGB1 => rgb_g_wire,
            CURREN => \N__35675\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__20028\,
            RGB0PWM => \N__47124\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18480\,
            in2 => \_gnd_net_\,
            in3 => \N__18733\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18471\,
            in2 => \N__18459\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18450\,
            in2 => \N__18438\,
            in3 => \N__18426\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18423\,
            in2 => \N__18411\,
            in3 => \N__18399\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18396\,
            in2 => \N__18384\,
            in3 => \N__18372\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18609\,
            in2 => \N__18758\,
            in3 => \N__18597\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18753\,
            in2 => \N__18594\,
            in3 => \N__18579\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18576\,
            in2 => \N__18759\,
            in3 => \N__18564\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18757\,
            in2 => \N__18561\,
            in3 => \N__18546\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18543\,
            in2 => \N__18734\,
            in3 => \N__18531\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18528\,
            in2 => \N__18738\,
            in3 => \N__18516\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18513\,
            in2 => \N__18735\,
            in3 => \N__18498\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18495\,
            in2 => \N__18739\,
            in3 => \N__18483\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18801\,
            in2 => \N__18736\,
            in3 => \N__18789\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18786\,
            in2 => \N__18740\,
            in3 => \N__18774\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18771\,
            in2 => \N__18737\,
            in3 => \N__18675\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18672\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20187\,
            in2 => \N__19454\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20155\,
            in2 => \N__18669\,
            in3 => \N__18654\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18651\,
            in2 => \N__21094\,
            in3 => \N__18642\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21022\,
            in2 => \N__18639\,
            in3 => \N__18627\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20942\,
            in2 => \N__18624\,
            in3 => \N__18942\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20862\,
            in2 => \N__18939\,
            in3 => \N__18927\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20795\,
            in2 => \N__18924\,
            in3 => \N__18909\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20727\,
            in2 => \N__18906\,
            in3 => \N__18891\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18888\,
            in2 => \N__20654\,
            in3 => \N__18876\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21529\,
            in2 => \N__18873\,
            in3 => \N__18858\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21477\,
            in2 => \N__18855\,
            in3 => \N__18837\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21436\,
            in2 => \N__18834\,
            in3 => \N__18819\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21370\,
            in2 => \N__18816\,
            in3 => \N__18804\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21308\,
            in2 => \N__19065\,
            in3 => \N__19053\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21247\,
            in2 => \N__19050\,
            in3 => \N__19038\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21195\,
            in2 => \N__19035\,
            in3 => \N__19020\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21141\,
            in2 => \N__19017\,
            in3 => \N__19002\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18999\,
            in2 => \N__21860\,
            in3 => \N__18990\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21804\,
            in2 => \N__18987\,
            in3 => \N__18975\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22773\,
            in2 => \N__18972\,
            in3 => \N__18960\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22744\,
            in2 => \N__18957\,
            in3 => \N__18945\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21768\,
            in2 => \N__19206\,
            in3 => \N__19194\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19191\,
            in2 => \N__21720\,
            in3 => \N__19182\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22815\,
            in2 => \N__19179\,
            in3 => \N__19164\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21639\,
            in2 => \N__19161\,
            in3 => \N__19146\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21591\,
            in2 => \N__19143\,
            in3 => \N__19131\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22110\,
            in2 => \N__19128\,
            in3 => \N__19113\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22071\,
            in2 => \N__19110\,
            in3 => \N__19098\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19095\,
            in2 => \N__22030\,
            in3 => \N__19086\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21982\,
            in2 => \N__19083\,
            in3 => \N__19068\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19284\,
            in1 => \N__22620\,
            in2 => \N__19275\,
            in3 => \N__19260\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001000"
        )
    port map (
            in0 => \N__20551\,
            in1 => \N__19257\,
            in2 => \N__20368\,
            in3 => \N__22652\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47516\,
            ce => 'H',
            sr => \N__47089\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111001000100"
        )
    port map (
            in0 => \N__20552\,
            in1 => \N__22650\,
            in2 => \N__20369\,
            in3 => \N__19251\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47516\,
            ce => 'H',
            sr => \N__47089\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22649\,
            in1 => \N__20555\,
            in2 => \N__19245\,
            in3 => \N__20315\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47516\,
            ce => 'H',
            sr => \N__47089\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__20553\,
            in1 => \N__22651\,
            in2 => \N__20370\,
            in3 => \N__19236\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47516\,
            ce => 'H',
            sr => \N__47089\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22648\,
            in1 => \N__20554\,
            in2 => \N__19227\,
            in3 => \N__20314\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47516\,
            ce => 'H',
            sr => \N__47089\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_1_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21251\,
            in1 => \N__21371\,
            in2 => \N__21551\,
            in3 => \N__22034\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19212\,
            in1 => \N__19551\,
            in2 => \N__19215\,
            in3 => \N__19314\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21209\,
            in1 => \N__21309\,
            in2 => \N__21441\,
            in3 => \N__21494\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21858\,
            in1 => \N__21817\,
            in2 => \N__21161\,
            in3 => \N__21773\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22664\,
            in1 => \N__21724\,
            in2 => \N__19317\,
            in3 => \N__19299\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21592\,
            in2 => \_gnd_net_\,
            in3 => \N__22737\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22076\,
            in1 => \N__22121\,
            in2 => \N__21651\,
            in3 => \N__21986\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22831\,
            in1 => \N__22786\,
            in2 => \N__19308\,
            in3 => \N__19305\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_1_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__26902\,
            in1 => \N__20995\,
            in2 => \_gnd_net_\,
            in3 => \N__19907\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20994\,
            in2 => \_gnd_net_\,
            in3 => \N__21064\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__19886\,
            in1 => \N__26903\,
            in2 => \N__19290\,
            in3 => \N__19677\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110010"
        )
    port map (
            in0 => \N__19343\,
            in1 => \N__19946\,
            in2 => \N__19287\,
            in3 => \N__21065\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19639\,
            in1 => \N__21951\,
            in2 => \N__19370\,
            in3 => \N__19330\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__47098\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010101000100"
        )
    port map (
            in0 => \N__26908\,
            in1 => \N__19960\,
            in2 => \N__19701\,
            in3 => \N__20931\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__47098\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19640\,
            in1 => \N__20583\,
            in2 => \N__19371\,
            in3 => \N__19331\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__47098\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__19329\,
            in1 => \N__20130\,
            in2 => \N__19363\,
            in3 => \N__19641\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__47098\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011111011"
        )
    port map (
            in0 => \N__21069\,
            in1 => \N__19344\,
            in2 => \N__19965\,
            in3 => \N__19332\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__47098\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__21003\,
            in1 => \N__19896\,
            in2 => \N__19702\,
            in3 => \N__19887\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47448\,
            ce => 'H',
            sr => \N__47098\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__26909\,
            in1 => \N__20844\,
            in2 => \N__19703\,
            in3 => \N__19963\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47442\,
            ce => 'H',
            sr => \N__47099\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19961\,
            in1 => \N__26910\,
            in2 => \N__20769\,
            in3 => \N__19699\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47442\,
            ce => 'H',
            sr => \N__47099\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000100"
        )
    port map (
            in0 => \N__26911\,
            in1 => \N__20691\,
            in2 => \N__19704\,
            in3 => \N__19964\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47442\,
            ce => 'H',
            sr => \N__47099\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000110010"
        )
    port map (
            in0 => \N__19962\,
            in1 => \N__26912\,
            in2 => \N__20622\,
            in3 => \N__19700\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47442\,
            ce => 'H',
            sr => \N__47099\
        );

    \rgb_drv_RNO_0_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__47123\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32673\,
            lcout => \N_38_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__20194\,
            in1 => \N__20523\,
            in2 => \N__19455\,
            in3 => \N__20378\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47547\,
            ce => 'H',
            sr => \N__47071\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22691\,
            in1 => \N__20520\,
            in2 => \N__19431\,
            in3 => \N__20375\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__20518\,
            in1 => \N__20371\,
            in2 => \_gnd_net_\,
            in3 => \N__19422\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__20516\,
            in1 => \N__22694\,
            in2 => \N__19416\,
            in3 => \N__20372\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22692\,
            in1 => \N__20521\,
            in2 => \N__19407\,
            in3 => \N__20376\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000010110001"
        )
    port map (
            in0 => \N__20519\,
            in1 => \N__22696\,
            in2 => \N__19398\,
            in3 => \N__20374\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__22693\,
            in1 => \N__20522\,
            in2 => \N__19389\,
            in3 => \N__20377\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__20517\,
            in1 => \N__22695\,
            in2 => \N__19380\,
            in3 => \N__20373\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47538\,
            ce => 'H',
            sr => \N__47074\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__22699\,
            in1 => \N__20514\,
            in2 => \N__20399\,
            in3 => \N__19539\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47529\,
            ce => 'H',
            sr => \N__47079\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__20512\,
            in1 => \N__22702\,
            in2 => \N__19533\,
            in3 => \N__20395\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47529\,
            ce => 'H',
            sr => \N__47079\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101010"
        )
    port map (
            in0 => \N__22700\,
            in1 => \N__19524\,
            in2 => \N__20400\,
            in3 => \N__20515\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47529\,
            ce => 'H',
            sr => \N__47079\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__20511\,
            in1 => \N__22701\,
            in2 => \N__19515\,
            in3 => \N__20394\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47529\,
            ce => 'H',
            sr => \N__47079\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__20513\,
            in1 => \N__22703\,
            in2 => \N__19506\,
            in3 => \N__20396\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47529\,
            ce => 'H',
            sr => \N__47079\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22655\,
            in1 => \N__20525\,
            in2 => \N__19494\,
            in3 => \N__20355\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001111100000"
        )
    port map (
            in0 => \N__20350\,
            in1 => \N__20557\,
            in2 => \N__19485\,
            in3 => \N__22660\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22656\,
            in1 => \N__20526\,
            in2 => \N__19476\,
            in3 => \N__20356\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20351\,
            in1 => \N__22657\,
            in2 => \N__20558\,
            in3 => \N__19467\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20352\,
            in1 => \N__22658\,
            in2 => \N__20559\,
            in3 => \N__19593\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22654\,
            in1 => \N__20524\,
            in2 => \N__19587\,
            in3 => \N__20354\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__20353\,
            in1 => \N__22659\,
            in2 => \N__20560\,
            in3 => \N__19578\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47517\,
            ce => 'H',
            sr => \N__47083\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__22653\,
            in1 => \N__20556\,
            in2 => \N__19572\,
            in3 => \N__20316\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47504\,
            ce => 'H',
            sr => \N__47087\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21300\,
            in2 => \_gnd_net_\,
            in3 => \N__21487\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21437\,
            in1 => \N__19608\,
            in2 => \N__19557\,
            in3 => \N__21981\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010111"
        )
    port map (
            in0 => \N__21106\,
            in1 => \N__20165\,
            in2 => \N__20209\,
            in3 => \N__21034\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__20647\,
            in2 => \N__19554\,
            in3 => \N__20878\,
            lcout => \current_shift_inst.PI_CTRL.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__20790\,
            in1 => \N__20956\,
            in2 => \_gnd_net_\,
            in3 => \N__20728\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20729\,
            in1 => \N__20791\,
            in2 => \N__20882\,
            in3 => \N__20646\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21107\,
            in1 => \N__21035\,
            in2 => \N__19629\,
            in3 => \N__20957\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21769\,
            in1 => \N__21859\,
            in2 => \N__21824\,
            in3 => \N__21160\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22026\,
            in1 => \N__21731\,
            in2 => \N__19626\,
            in3 => \N__19623\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19617\,
            in1 => \N__22554\,
            in2 => \N__19611\,
            in3 => \N__19602\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21243\,
            in1 => \N__21360\,
            in2 => \N__21210\,
            in3 => \N__21535\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22117\,
            in1 => \N__21643\,
            in2 => \N__21608\,
            in3 => \N__22072\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21326\,
            in1 => \N__21668\,
            in2 => \N__21687\,
            in3 => \N__21272\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__20608\,
            in1 => \_gnd_net_\,
            in2 => \N__20926\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__20683\,
            in1 => \N__20764\,
            in2 => \N__19596\,
            in3 => \N__20833\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21398\,
            in2 => \_gnd_net_\,
            in3 => \N__21887\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21458\,
            in1 => \N__22326\,
            in2 => \N__19728\,
            in3 => \N__19725\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21273\,
            in1 => \N__21935\,
            in2 => \N__21330\,
            in3 => \N__21920\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21669\,
            in1 => \N__21683\,
            in2 => \N__22343\,
            in3 => \N__21902\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22242\,
            in1 => \N__19719\,
            in2 => \N__19713\,
            in3 => \N__22371\,
            lcout => \current_shift_inst.PI_CTRL.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22404\,
            in2 => \_gnd_net_\,
            in3 => \N__22389\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21459\,
            in1 => \N__21402\,
            in2 => \N__19656\,
            in3 => \N__21870\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21909\,
            in1 => \N__19653\,
            in2 => \N__19644\,
            in3 => \N__22308\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19913\,
            in2 => \N__26904\,
            in3 => \N__19945\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__21002\,
            in1 => \N__19947\,
            in2 => \N__19917\,
            in3 => \N__26886\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20687\,
            in2 => \_gnd_net_\,
            in3 => \N__20927\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20765\,
            in1 => \N__20840\,
            in2 => \N__19890\,
            in3 => \N__20615\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19871\,
            in1 => \N__19856\,
            in2 => \_gnd_net_\,
            in3 => \N__19838\,
            lcout => \pwm_generator_inst.un1_duty_inputlt3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19753\,
            in1 => \N__19823\,
            in2 => \N__19784\,
            in3 => \N__19801\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19822\,
            in2 => \_gnd_net_\,
            in3 => \N__20047\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__19802\,
            in1 => \N__19780\,
            in2 => \N__19761\,
            in3 => \N__19754\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111011"
        )
    port map (
            in0 => \N__19737\,
            in1 => \N__20074\,
            in2 => \N__19731\,
            in3 => \N__20101\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__20112\,
            in1 => \N__20106\,
            in2 => \N__20082\,
            in3 => \N__20054\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rgb_drv_RNO_LC_2_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__47122\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32672\,
            lcout => \rgb_drv_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20019\,
            in1 => \N__20568\,
            in2 => \_gnd_net_\,
            in3 => \N__20397\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47539\,
            ce => 'H',
            sr => \N__47067\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011010001"
        )
    port map (
            in0 => \N__22704\,
            in1 => \N__20561\,
            in2 => \N__20010\,
            in3 => \N__20398\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47530\,
            ce => 'H',
            sr => \N__47072\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__20386\,
            in1 => \N__22705\,
            in2 => \N__19995\,
            in3 => \N__20565\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47518\,
            ce => 'H',
            sr => \N__47075\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22538\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47505\,
            ce => 'H',
            sr => \N__47080\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23027\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47505\,
            ce => 'H',
            sr => \N__47080\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22698\,
            in1 => \N__20567\,
            in2 => \N__19980\,
            in3 => \N__20385\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47505\,
            ce => 'H',
            sr => \N__47080\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22490\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47505\,
            ce => 'H',
            sr => \N__47080\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_3_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22433\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22949\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22922\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__20228\,
            in1 => \N__20213\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22467\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22871\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23003\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011100010"
        )
    port map (
            in0 => \N__22706\,
            in1 => \N__20566\,
            in2 => \N__20415\,
            in3 => \N__20387\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47492\,
            ce => 'H',
            sr => \N__47084\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20229\,
            in2 => \N__20214\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22236\,
            in2 => \N__20166\,
            in3 => \N__20115\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21117\,
            in2 => \N__21108\,
            in3 => \N__21045\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21042\,
            in2 => \N__21036\,
            in3 => \N__20973\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20970\,
            in2 => \N__20964\,
            in3 => \N__20895\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20892\,
            in2 => \N__20883\,
            in3 => \N__20811\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20808\,
            in2 => \N__20802\,
            in3 => \N__20733\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22839\,
            in2 => \N__20730\,
            in3 => \N__20658\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__47478\,
            ce => 'H',
            sr => \N__47088\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23046\,
            in2 => \N__20655\,
            in3 => \N__20586\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21561\,
            in2 => \N__21552\,
            in3 => \N__21510\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21507\,
            in2 => \N__21498\,
            in3 => \N__21444\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21435\,
            in2 => \N__22134\,
            in3 => \N__21384\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21381\,
            in2 => \N__21372\,
            in3 => \N__21312\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21301\,
            in2 => \N__22193\,
            in3 => \N__21258\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22157\,
            in2 => \N__21255\,
            in3 => \N__21213\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21208\,
            in2 => \N__22194\,
            in3 => \N__21168\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__47466\,
            ce => 'H',
            sr => \N__47090\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22195\,
            in2 => \N__21165\,
            in3 => \N__21120\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21864\,
            in2 => \N__22224\,
            in3 => \N__21828\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22199\,
            in2 => \N__21825\,
            in3 => \N__21783\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22791\,
            in2 => \N__22225\,
            in3 => \N__21780\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22203\,
            in2 => \N__22751\,
            in3 => \N__21777\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21774\,
            in2 => \N__22226\,
            in3 => \N__21735\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22207\,
            in2 => \N__21732\,
            in3 => \N__21672\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22833\,
            in2 => \N__22227\,
            in3 => \N__21654\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__47458\,
            ce => 'H',
            sr => \N__47093\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21650\,
            in2 => \N__22228\,
            in3 => \N__21612\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22214\,
            in2 => \N__21609\,
            in3 => \N__21564\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22122\,
            in2 => \N__22229\,
            in3 => \N__22083\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22218\,
            in2 => \N__22080\,
            in3 => \N__22038\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22035\,
            in2 => \N__22230\,
            in3 => \N__21996\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22222\,
            in2 => \N__21993\,
            in3 => \N__21957\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__22223\,
            in1 => \N__22707\,
            in2 => \_gnd_net_\,
            in3 => \N__21954\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22848\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47449\,
            ce => 'H',
            sr => \N__47094\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22251\,
            in1 => \N__21939\,
            in2 => \N__22266\,
            in3 => \N__21924\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22290\,
            in1 => \N__21903\,
            in2 => \N__21891\,
            in3 => \N__22302\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22353\,
            in1 => \N__22403\,
            in2 => \N__22365\,
            in3 => \N__22388\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22364\,
            in2 => \_gnd_net_\,
            in3 => \N__22352\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22344\,
            in1 => \N__22325\,
            in2 => \N__22311\,
            in3 => \N__22278\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22301\,
            in1 => \N__22289\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22277\,
            in1 => \N__22262\,
            in2 => \N__22254\,
            in3 => \N__22250\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22511\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47479\,
            ce => 'H',
            sr => \N__47081\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23091\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47479\,
            ce => 'H',
            sr => \N__47081\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22892\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47479\,
            ce => 'H',
            sr => \N__47081\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24380\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => 'H',
            sr => \N__47085\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22973\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47467\,
            ce => 'H',
            sr => \N__47085\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22832\,
            in1 => \N__22790\,
            in2 => \N__22752\,
            in3 => \N__22697\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22545\,
            in2 => \_gnd_net_\,
            in3 => \N__24114\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24105\,
            in2 => \_gnd_net_\,
            in3 => \N__22521\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24348\,
            in2 => \_gnd_net_\,
            in3 => \N__22497\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24336\,
            in2 => \_gnd_net_\,
            in3 => \N__22470\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24324\,
            in2 => \_gnd_net_\,
            in3 => \N__22437\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24312\,
            in2 => \_gnd_net_\,
            in3 => \N__22407\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24300\,
            in2 => \_gnd_net_\,
            in3 => \N__23007\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24288\,
            in2 => \_gnd_net_\,
            in3 => \N__22980\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__47480\,
            ce => 'H',
            sr => \N__47073\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24276\,
            in2 => \_gnd_net_\,
            in3 => \N__22959\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24264\,
            in2 => \_gnd_net_\,
            in3 => \N__22956\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24447\,
            in2 => \_gnd_net_\,
            in3 => \N__22929\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24435\,
            in2 => \_gnd_net_\,
            in3 => \N__22902\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24423\,
            in2 => \_gnd_net_\,
            in3 => \N__22878\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23352\,
            in2 => \_gnd_net_\,
            in3 => \N__22851\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24408\,
            in2 => \_gnd_net_\,
            in3 => \N__23163\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47468\,
            ce => 'H',
            sr => \N__47076\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23066\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47450\,
            ce => 'H',
            sr => \N__47086\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26514\,
            in1 => \N__26539\,
            in2 => \_gnd_net_\,
            in3 => \N__41184\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47548\,
            ce => \N__32100\,
            sr => \N__47029\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41133\,
            in1 => \N__24961\,
            in2 => \_gnd_net_\,
            in3 => \N__24940\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47540\,
            ce => \N__32112\,
            sr => \N__47035\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25093\,
            in1 => \N__25068\,
            in2 => \_gnd_net_\,
            in3 => \N__41132\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25015\,
            in1 => \N__24980\,
            in2 => \_gnd_net_\,
            in3 => \N__41181\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => \elapsed_time_ns_1_RNI02CN9_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41182\,
            in1 => \_gnd_net_\,
            in2 => \N__23037\,
            in3 => \N__25016\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47531\,
            ce => \N__32101\,
            sr => \N__47041\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23653\,
            in2 => \N__23703\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23632\,
            in2 => \N__23679\,
            in3 => \N__23034\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23654\,
            in2 => \N__23612\,
            in3 => \N__23193\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23584\,
            in2 => \N__23637\,
            in3 => \N__23190\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23563\,
            in2 => \N__23613\,
            in3 => \N__23187\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23887\,
            in2 => \N__23589\,
            in3 => \N__23184\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23564\,
            in2 => \N__23871\,
            in3 => \N__23181\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23888\,
            in2 => \N__23841\,
            in3 => \N__23178\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47519\,
            ce => \N__25221\,
            sr => \N__47046\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23809\,
            in2 => \N__23870\,
            in3 => \N__23175\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23788\,
            in2 => \N__23840\,
            in3 => \N__23172\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23810\,
            in2 => \N__23768\,
            in3 => \N__23169\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23740\,
            in2 => \N__23793\,
            in3 => \N__23166\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23719\,
            in2 => \N__23769\,
            in3 => \N__23220\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24091\,
            in2 => \N__23745\,
            in3 => \N__23217\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23720\,
            in2 => \N__24075\,
            in3 => \N__23214\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24092\,
            in2 => \N__24045\,
            in3 => \N__23211\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47506\,
            ce => \N__25220\,
            sr => \N__47052\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24013\,
            in2 => \N__24074\,
            in3 => \N__23208\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23992\,
            in2 => \N__24044\,
            in3 => \N__23205\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24014\,
            in2 => \N__23972\,
            in3 => \N__23202\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23944\,
            in2 => \N__23997\,
            in3 => \N__23199\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23923\,
            in2 => \N__23973\,
            in3 => \N__23196\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23905\,
            in2 => \N__23949\,
            in3 => \N__23244\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23924\,
            in2 => \N__24252\,
            in3 => \N__23241\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23906\,
            in2 => \N__24222\,
            in3 => \N__23238\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47493\,
            ce => \N__25218\,
            sr => \N__47056\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24187\,
            in2 => \N__24251\,
            in3 => \N__23235\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47481\,
            ce => \N__25217\,
            sr => \N__47059\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24163\,
            in2 => \N__24221\,
            in3 => \N__23232\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47481\,
            ce => \N__25217\,
            sr => \N__47059\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24143\,
            in2 => \N__24192\,
            in3 => \N__23229\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47481\,
            ce => \N__25217\,
            sr => \N__47059\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24125\,
            in2 => \N__24168\,
            in3 => \N__23226\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47481\,
            ce => \N__25217\,
            sr => \N__47059\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23223\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47481\,
            ce => \N__25217\,
            sr => \N__47059\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25906\,
            in1 => \N__25867\,
            in2 => \_gnd_net_\,
            in3 => \N__41169\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25395\,
            in1 => \N__41196\,
            in2 => \_gnd_net_\,
            in3 => \N__25416\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47451\,
            ce => \N__32111\,
            sr => \N__47068\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24404\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42407\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_7_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__27307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27269\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23328\,
            in3 => \N__23343\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23307\,
            in2 => \_gnd_net_\,
            in3 => \N__23319\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23286\,
            in2 => \_gnd_net_\,
            in3 => \N__23301\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23265\,
            in2 => \_gnd_net_\,
            in3 => \N__23280\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23469\,
            in2 => \_gnd_net_\,
            in3 => \N__23259\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23448\,
            in2 => \_gnd_net_\,
            in3 => \N__23463\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23427\,
            in2 => \_gnd_net_\,
            in3 => \N__23442\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23406\,
            in2 => \_gnd_net_\,
            in3 => \N__23421\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23385\,
            in2 => \_gnd_net_\,
            in3 => \N__23400\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23379\,
            in1 => \N__23367\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_7_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27308\,
            in2 => \_gnd_net_\,
            in3 => \N__23361\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_7_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__29873\,
            in1 => \N__25649\,
            in2 => \_gnd_net_\,
            in3 => \N__23358\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_7_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29932\,
            in2 => \_gnd_net_\,
            in3 => \N__23355\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_7_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27226\,
            in2 => \_gnd_net_\,
            in3 => \N__23499\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_7_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27325\,
            in2 => \_gnd_net_\,
            in3 => \N__23496\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_7_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29776\,
            in2 => \_gnd_net_\,
            in3 => \N__23493\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_7_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27388\,
            in2 => \_gnd_net_\,
            in3 => \N__23490\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_7_28_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27427\,
            in2 => \_gnd_net_\,
            in3 => \N__23487\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25699\,
            in2 => \_gnd_net_\,
            in3 => \N__23484\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23481\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23478\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47552\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__28295\,
            in1 => \N__23523\,
            in2 => \N__28323\,
            in3 => \N__23511\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__23510\,
            in1 => \N__28322\,
            in2 => \N__28299\,
            in3 => \N__23522\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26624\,
            in1 => \N__26590\,
            in2 => \_gnd_net_\,
            in3 => \N__41138\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47541\,
            ce => \N__32106\,
            sr => \N__47023\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26170\,
            in1 => \N__26217\,
            in2 => \N__25071\,
            in3 => \N__26286\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23547\,
            in1 => \N__23535\,
            in2 => \N__23502\,
            in3 => \N__23529\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25384\,
            in2 => \_gnd_net_\,
            in3 => \N__26046\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24965\,
            in1 => \N__24939\,
            in2 => \_gnd_net_\,
            in3 => \N__41135\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__24612\,
            in1 => \N__26355\,
            in2 => \_gnd_net_\,
            in3 => \N__23541\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24581\,
            in1 => \N__24613\,
            in2 => \_gnd_net_\,
            in3 => \N__41136\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41134\,
            in1 => \N__26543\,
            in2 => \_gnd_net_\,
            in3 => \N__26521\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26805\,
            in1 => \N__24768\,
            in2 => \N__27080\,
            in3 => \N__41235\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25126\,
            in1 => \N__26103\,
            in2 => \N__24529\,
            in3 => \N__24840\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__24722\,
            in1 => \_gnd_net_\,
            in2 => \N__41187\,
            in3 => \N__24697\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24522\,
            in1 => \N__41143\,
            in2 => \_gnd_net_\,
            in3 => \N__24560\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25866\,
            in1 => \N__26748\,
            in2 => \N__26523\,
            in3 => \N__26580\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26806\,
            in1 => \N__41142\,
            in2 => \_gnd_net_\,
            in3 => \N__26831\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24873\,
            in1 => \N__24696\,
            in2 => \N__24944\,
            in3 => \N__25011\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47507\,
            ce => \N__25219\,
            sr => \N__47042\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23678\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47507\,
            ce => \N__25219\,
            sr => \N__47042\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24818\,
            in1 => \N__24841\,
            in2 => \_gnd_net_\,
            in3 => \N__41160\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41159\,
            in1 => \N__26080\,
            in2 => \_gnd_net_\,
            in3 => \N__26104\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25163\,
            in1 => \N__25127\,
            in2 => \_gnd_net_\,
            in3 => \N__41161\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25324\,
            in1 => \N__23698\,
            in2 => \_gnd_net_\,
            in3 => \N__23682\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25347\,
            in1 => \N__23674\,
            in2 => \_gnd_net_\,
            in3 => \N__23658\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25325\,
            in1 => \N__23655\,
            in2 => \_gnd_net_\,
            in3 => \N__23640\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25348\,
            in1 => \N__23633\,
            in2 => \_gnd_net_\,
            in3 => \N__23616\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25326\,
            in1 => \N__23611\,
            in2 => \_gnd_net_\,
            in3 => \N__23592\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25349\,
            in1 => \N__23585\,
            in2 => \_gnd_net_\,
            in3 => \N__23568\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25327\,
            in1 => \N__23565\,
            in2 => \_gnd_net_\,
            in3 => \N__23550\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25350\,
            in1 => \N__23889\,
            in2 => \_gnd_net_\,
            in3 => \N__23874\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__47494\,
            ce => \N__25548\,
            sr => \N__47047\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25323\,
            in1 => \N__23863\,
            in2 => \_gnd_net_\,
            in3 => \N__23844\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25331\,
            in1 => \N__23833\,
            in2 => \_gnd_net_\,
            in3 => \N__23814\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25320\,
            in1 => \N__23811\,
            in2 => \_gnd_net_\,
            in3 => \N__23796\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25328\,
            in1 => \N__23789\,
            in2 => \_gnd_net_\,
            in3 => \N__23772\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25321\,
            in1 => \N__23767\,
            in2 => \_gnd_net_\,
            in3 => \N__23748\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25329\,
            in1 => \N__23741\,
            in2 => \_gnd_net_\,
            in3 => \N__23724\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25322\,
            in1 => \N__23721\,
            in2 => \_gnd_net_\,
            in3 => \N__23706\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25330\,
            in1 => \N__24093\,
            in2 => \_gnd_net_\,
            in3 => \N__24078\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__47482\,
            ce => \N__25547\,
            sr => \N__47053\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25316\,
            in1 => \N__24067\,
            in2 => \_gnd_net_\,
            in3 => \N__24048\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25334\,
            in1 => \N__24037\,
            in2 => \_gnd_net_\,
            in3 => \N__24018\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25317\,
            in1 => \N__24015\,
            in2 => \_gnd_net_\,
            in3 => \N__24000\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25335\,
            in1 => \N__23993\,
            in2 => \_gnd_net_\,
            in3 => \N__23976\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25318\,
            in1 => \N__23971\,
            in2 => \_gnd_net_\,
            in3 => \N__23952\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25336\,
            in1 => \N__23945\,
            in2 => \_gnd_net_\,
            in3 => \N__23928\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25319\,
            in1 => \N__23925\,
            in2 => \_gnd_net_\,
            in3 => \N__23910\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25337\,
            in1 => \N__23907\,
            in2 => \_gnd_net_\,
            in3 => \N__23892\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__47469\,
            ce => \N__25546\,
            sr => \N__47057\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25312\,
            in1 => \N__24244\,
            in2 => \_gnd_net_\,
            in3 => \N__24225\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__47459\,
            ce => \N__25536\,
            sr => \N__47060\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25332\,
            in1 => \N__24214\,
            in2 => \_gnd_net_\,
            in3 => \N__24195\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__47459\,
            ce => \N__25536\,
            sr => \N__47060\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25313\,
            in1 => \N__24188\,
            in2 => \_gnd_net_\,
            in3 => \N__24171\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__47459\,
            ce => \N__25536\,
            sr => \N__47060\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25333\,
            in1 => \N__24164\,
            in2 => \_gnd_net_\,
            in3 => \N__24147\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__47459\,
            ce => \N__25536\,
            sr => \N__47060\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25314\,
            in1 => \N__24144\,
            in2 => \_gnd_net_\,
            in3 => \N__24132\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__47459\,
            ce => \N__25536\,
            sr => \N__47060\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__24126\,
            in1 => \N__25315\,
            in2 => \_gnd_net_\,
            in3 => \N__24129\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47459\,
            ce => \N__25536\,
            sr => \N__47060\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25496\,
            in2 => \N__25473\,
            in3 => \N__25471\,
            lcout => \current_shift_inst.control_input_18\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25503\,
            in2 => \_gnd_net_\,
            in3 => \N__24096\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25485\,
            in2 => \_gnd_net_\,
            in3 => \N__24339\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25479\,
            in2 => \_gnd_net_\,
            in3 => \N__24327\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29418\,
            in2 => \_gnd_net_\,
            in3 => \N__24315\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25452\,
            in2 => \_gnd_net_\,
            in3 => \N__24303\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29439\,
            in2 => \_gnd_net_\,
            in3 => \N__24291\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25446\,
            in2 => \_gnd_net_\,
            in3 => \N__24279\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26949\,
            in2 => \_gnd_net_\,
            in3 => \N__24267\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26937\,
            in2 => \_gnd_net_\,
            in3 => \N__24255\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26925\,
            in2 => \_gnd_net_\,
            in3 => \N__24438\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29457\,
            in2 => \_gnd_net_\,
            in3 => \N__24426\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24393\,
            in2 => \_gnd_net_\,
            in3 => \N__24414\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35298\,
            in2 => \_gnd_net_\,
            in3 => \N__24411\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35297\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25497\,
            in2 => \_gnd_net_\,
            in3 => \N__25472\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47437\,
            ce => 'H',
            sr => \N__47069\
        );

    \phase_controller_inst2.S2_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41955\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47424\,
            ce => 'H',
            sr => \N__47091\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_8_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__27329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27344\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_8_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__27230\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27248\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_8_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__29780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29753\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_8_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27392\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_8_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29906\,
            in2 => \_gnd_net_\,
            in3 => \N__29936\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_8_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27446\,
            in2 => \_gnd_net_\,
            in3 => \N__27431\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_8_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__25700\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25712\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_8_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47559\,
            lcout => \GB_BUFFER_clock_output_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27097\,
            in1 => \N__27079\,
            in2 => \_gnd_net_\,
            in3 => \N__41183\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47553\,
            ce => \N__32071\,
            sr => \N__46996\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24797\,
            in1 => \N__24776\,
            in2 => \_gnd_net_\,
            in3 => \N__41137\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41109\,
            in1 => \N__24793\,
            in2 => \_gnd_net_\,
            in3 => \N__24777\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47542\,
            ce => \N__32018\,
            sr => \N__47010\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26763\,
            in1 => \N__26717\,
            in2 => \_gnd_net_\,
            in3 => \N__41110\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47542\,
            ce => \N__32018\,
            sr => \N__47010\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__28430\,
            in1 => \N__28406\,
            in2 => \N__24498\,
            in3 => \N__24486\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40949\,
            in1 => \N__24905\,
            in2 => \_gnd_net_\,
            in3 => \N__24883\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__24485\,
            in1 => \N__28431\,
            in2 => \N__28410\,
            in3 => \N__24494\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26177\,
            in1 => \N__26138\,
            in2 => \_gnd_net_\,
            in3 => \N__40950\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => \elapsed_time_ns_1_RNI68CN9_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__40951\,
            in1 => \_gnd_net_\,
            in2 => \N__24501\,
            in3 => \N__26178\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47532\,
            ce => \N__32105\,
            sr => \N__47016\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24621\,
            in1 => \N__24577\,
            in2 => \_gnd_net_\,
            in3 => \N__40993\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47520\,
            ce => \N__32107\,
            sr => \N__47024\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40991\,
            in1 => \N__26239\,
            in2 => \_gnd_net_\,
            in3 => \N__26222\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47520\,
            ce => \N__32107\,
            sr => \N__47024\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40992\,
            in2 => \N__26685\,
            in3 => \N__26661\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47520\,
            ce => \N__32107\,
            sr => \N__47024\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26827\,
            in1 => \N__26811\,
            in2 => \_gnd_net_\,
            in3 => \N__40994\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47520\,
            ce => \N__32107\,
            sr => \N__47024\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40990\,
            in1 => \N__24901\,
            in2 => \_gnd_net_\,
            in3 => \N__24885\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47520\,
            ce => \N__32107\,
            sr => \N__47024\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25787\,
            in1 => \N__25981\,
            in2 => \_gnd_net_\,
            in3 => \N__40995\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47520\,
            ce => \N__32107\,
            sr => \N__47024\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40996\,
            in1 => \N__24814\,
            in2 => \_gnd_net_\,
            in3 => \N__24842\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47508\,
            ce => \N__32079\,
            sr => \N__47030\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24637\,
            in1 => \N__24668\,
            in2 => \_gnd_net_\,
            in3 => \N__40999\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47508\,
            ce => \N__32079\,
            sr => \N__47030\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40998\,
            in1 => \N__24556\,
            in2 => \_gnd_net_\,
            in3 => \N__24540\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47508\,
            ce => \N__32079\,
            sr => \N__47030\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24718\,
            in1 => \N__24702\,
            in2 => \_gnd_net_\,
            in3 => \N__41000\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47508\,
            ce => \N__32079\,
            sr => \N__47030\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40997\,
            in1 => \N__25159\,
            in2 => \_gnd_net_\,
            in3 => \N__25139\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47508\,
            ce => \N__32079\,
            sr => \N__47030\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25100\,
            in1 => \N__25070\,
            in2 => \_gnd_net_\,
            in3 => \N__41001\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47508\,
            ce => \N__32079\,
            sr => \N__47030\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26424\,
            in1 => \N__26390\,
            in2 => \N__26664\,
            in3 => \N__24660\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24639\,
            in1 => \N__24661\,
            in2 => \_gnd_net_\,
            in3 => \N__41162\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26425\,
            in1 => \N__26459\,
            in2 => \_gnd_net_\,
            in3 => \N__41163\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47495\,
            ce => \N__32070\,
            sr => \N__47036\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26391\,
            in1 => \N__41167\,
            in2 => \_gnd_net_\,
            in3 => \N__26406\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47495\,
            ce => \N__32070\,
            sr => \N__47036\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24798\,
            in1 => \N__24772\,
            in2 => \_gnd_net_\,
            in3 => \N__41127\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41121\,
            in1 => \N__24726\,
            in2 => \_gnd_net_\,
            in3 => \N__24701\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24669\,
            in1 => \N__24638\,
            in2 => \_gnd_net_\,
            in3 => \N__41125\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41122\,
            in1 => \N__24620\,
            in2 => \_gnd_net_\,
            in3 => \N__24582\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25907\,
            in1 => \N__25874\,
            in2 => \_gnd_net_\,
            in3 => \N__41126\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41124\,
            in1 => \N__26013\,
            in2 => \_gnd_net_\,
            in3 => \N__26057\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24561\,
            in1 => \N__24536\,
            in2 => \_gnd_net_\,
            in3 => \N__41128\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41123\,
            in1 => \N__25164\,
            in2 => \_gnd_net_\,
            in3 => \N__25143\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47483\,
            ce => \N__27019\,
            sr => \N__47043\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__31089\,
            in1 => \N__25110\,
            in2 => \N__25029\,
            in3 => \N__31112\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__25109\,
            in1 => \N__31088\,
            in2 => \N__31116\,
            in3 => \N__25025\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__41179\,
            in2 => \_gnd_net_\,
            in3 => \N__25069\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__27017\,
            sr => \N__47048\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25017\,
            in1 => \N__24987\,
            in2 => \_gnd_net_\,
            in3 => \N__41165\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__27017\,
            sr => \N__47048\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41164\,
            in1 => \N__24969\,
            in2 => \_gnd_net_\,
            in3 => \N__24945\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__27017\,
            sr => \N__47048\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24906\,
            in1 => \N__24884\,
            in2 => \_gnd_net_\,
            in3 => \N__41166\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__27017\,
            sr => \N__47048\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24846\,
            in1 => \N__41180\,
            in2 => \_gnd_net_\,
            in3 => \N__24819\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47470\,
            ce => \N__27017\,
            sr => \N__47048\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__31016\,
            in1 => \N__30989\,
            in2 => \N__25440\,
            in3 => \N__25425\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__25424\,
            in1 => \N__31017\,
            in2 => \N__30993\,
            in3 => \N__25436\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41190\,
            in1 => \N__26289\,
            in2 => \_gnd_net_\,
            in3 => \N__25833\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__27015\,
            sr => \N__47054\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41191\,
            in1 => \N__25982\,
            in2 => \_gnd_net_\,
            in3 => \N__25794\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__27015\,
            sr => \N__47054\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25393\,
            in1 => \N__41189\,
            in2 => \_gnd_net_\,
            in3 => \N__25409\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => \elapsed_time_ns_1_RNIK63T9_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41192\,
            in1 => \_gnd_net_\,
            in2 => \N__25398\,
            in3 => \N__25394\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47460\,
            ce => \N__27015\,
            sr => \N__47054\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25362\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41170\,
            in1 => \N__26356\,
            in2 => \_gnd_net_\,
            in3 => \N__26311\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26964\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26966\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28142\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_198_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26965\,
            in2 => \N__28146\,
            in3 => \N__29732\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_199_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26458\,
            in1 => \N__26436\,
            in2 => \_gnd_net_\,
            in3 => \N__41188\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__35286\,
            in1 => \N__31578\,
            in2 => \_gnd_net_\,
            in3 => \N__29367\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31593\,
            in1 => \N__29256\,
            in2 => \_gnd_net_\,
            in3 => \N__35284\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__35287\,
            in1 => \N__31563\,
            in2 => \_gnd_net_\,
            in3 => \N__29352\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31548\,
            in1 => \N__29337\,
            in2 => \_gnd_net_\,
            in3 => \N__35288\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35285\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.N_1288_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31680\,
            in1 => \N__29319\,
            in2 => \_gnd_net_\,
            in3 => \N__35289\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31653\,
            in1 => \N__29301\,
            in2 => \_gnd_net_\,
            in3 => \N__35290\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25650\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25617\,
            in2 => \_gnd_net_\,
            in3 => \N__25602\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25599\,
            in2 => \_gnd_net_\,
            in3 => \N__25584\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25581\,
            in2 => \_gnd_net_\,
            in3 => \N__25566\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27159\,
            in2 => \_gnd_net_\,
            in3 => \N__25563\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35467\,
            in2 => \N__27114\,
            in3 => \N__25560\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27798\,
            in2 => \N__35538\,
            in3 => \N__25557\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35471\,
            in2 => \N__27753\,
            in3 => \N__25554\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27699\,
            in2 => \_gnd_net_\,
            in3 => \N__25551\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27651\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27606\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27567\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27522\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28071\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28041\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28014\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27984\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27954\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27924\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27858\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25719\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__25716\,
            in1 => \N__29831\,
            in2 => \N__25701\,
            in3 => \N__25680\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100010000"
        )
    port map (
            in0 => \N__28272\,
            in1 => \N__28250\,
            in2 => \N__25662\,
            in3 => \N__25671\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101111"
        )
    port map (
            in0 => \N__25670\,
            in1 => \N__25658\,
            in2 => \N__28251\,
            in3 => \N__28271\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__27101\,
            in1 => \N__27081\,
            in2 => \_gnd_net_\,
            in3 => \N__41092\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41093\,
            in1 => \N__29681\,
            in2 => \_gnd_net_\,
            in3 => \N__29635\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000010"
        )
    port map (
            in0 => \N__25812\,
            in1 => \N__28226\,
            in2 => \N__28562\,
            in3 => \N__25803\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26364\,
            in1 => \N__26319\,
            in2 => \_gnd_net_\,
            in3 => \N__41105\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47521\,
            ce => \N__32049\,
            sr => \N__46997\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__25811\,
            in1 => \N__28227\,
            in2 => \N__28563\,
            in3 => \N__25802\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25786\,
            in1 => \N__25983\,
            in2 => \_gnd_net_\,
            in3 => \N__41104\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__25755\,
            in1 => \N__28531\,
            in2 => \N__25767\,
            in3 => \N__28513\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101001101"
        )
    port map (
            in0 => \N__28532\,
            in1 => \N__25766\,
            in2 => \N__28515\,
            in3 => \N__25754\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26008\,
            in1 => \N__26058\,
            in2 => \_gnd_net_\,
            in3 => \N__41002\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47510\,
            ce => \N__32080\,
            sr => \N__47005\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26623\,
            in1 => \N__26595\,
            in2 => \_gnd_net_\,
            in3 => \N__40946\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101110001"
        )
    port map (
            in0 => \N__28187\,
            in1 => \N__28165\,
            in2 => \N__25746\,
            in3 => \N__25730\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001110"
        )
    port map (
            in0 => \N__25745\,
            in1 => \N__25731\,
            in2 => \N__28167\,
            in3 => \N__28188\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40947\,
            in1 => \N__26243\,
            in2 => \_gnd_net_\,
            in3 => \N__26218\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26012\,
            in1 => \N__26056\,
            in2 => \_gnd_net_\,
            in3 => \N__40948\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25992\,
            in1 => \N__25977\,
            in2 => \N__29680\,
            in3 => \N__25944\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__28477\,
            in1 => \N__25935\,
            in2 => \N__25926\,
            in3 => \N__25923\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26758\,
            in2 => \N__25914\,
            in3 => \N__26716\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__26253\,
            in1 => \N__25841\,
            in2 => \N__28385\,
            in3 => \N__28352\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011101111"
        )
    port map (
            in0 => \N__25842\,
            in1 => \N__26252\,
            in2 => \N__28386\,
            in3 => \N__28353\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40957\,
            in1 => \N__25911\,
            in2 => \_gnd_net_\,
            in3 => \N__25878\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47484\,
            ce => \N__32078\,
            sr => \N__47017\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26287\,
            in1 => \N__40955\,
            in2 => \_gnd_net_\,
            in3 => \N__25826\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__40956\,
            in1 => \_gnd_net_\,
            in2 => \N__25815\,
            in3 => \N__26288\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47484\,
            ce => \N__32078\,
            sr => \N__47017\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26115\,
            in1 => \_gnd_net_\,
            in2 => \N__41111\,
            in3 => \N__26085\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47484\,
            ce => \N__32078\,
            sr => \N__47017\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__31067\,
            in1 => \N__31040\,
            in2 => \N__26127\,
            in3 => \N__26187\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__26186\,
            in1 => \N__31068\,
            in2 => \N__31044\,
            in3 => \N__26123\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26244\,
            in1 => \N__26223\,
            in2 => \_gnd_net_\,
            in3 => \N__41119\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47471\,
            ce => \N__27021\,
            sr => \N__47025\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41115\,
            in1 => \N__26176\,
            in2 => \_gnd_net_\,
            in3 => \N__26142\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47471\,
            ce => \N__27021\,
            sr => \N__47025\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26114\,
            in1 => \N__26081\,
            in2 => \_gnd_net_\,
            in3 => \N__41120\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47471\,
            ce => \N__27021\,
            sr => \N__47025\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29676\,
            in2 => \N__41185\,
            in3 => \N__29637\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47471\,
            ce => \N__27021\,
            sr => \N__47025\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__31347\,
            in1 => \N__31370\,
            in2 => \N__26475\,
            in3 => \N__26556\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26555\,
            in1 => \N__31346\,
            in2 => \N__31374\,
            in3 => \N__26471\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41096\,
            in1 => \N__26625\,
            in2 => \_gnd_net_\,
            in3 => \N__26594\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47461\,
            ce => \N__27020\,
            sr => \N__47031\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26547\,
            in1 => \N__26522\,
            in2 => \_gnd_net_\,
            in3 => \N__41098\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47461\,
            ce => \N__27020\,
            sr => \N__47031\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41097\,
            in1 => \N__26463\,
            in2 => \_gnd_net_\,
            in3 => \N__26435\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47461\,
            ce => \N__27020\,
            sr => \N__47031\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26388\,
            in1 => \N__26405\,
            in2 => \_gnd_net_\,
            in3 => \N__41094\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => \elapsed_time_ns_1_RNIUVBN9_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__41095\,
            in1 => \_gnd_net_\,
            in2 => \N__26394\,
            in3 => \N__26389\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47461\,
            ce => \N__27020\,
            sr => \N__47031\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__26993\,
            in1 => \N__26979\,
            in2 => \N__31245\,
            in3 => \N__31275\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41175\,
            in1 => \N__26363\,
            in2 => \_gnd_net_\,
            in3 => \N__26312\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__27018\,
            sr => \N__47037\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26843\,
            in1 => \N__31184\,
            in2 => \N__31212\,
            in3 => \N__26771\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__31185\,
            in1 => \N__31208\,
            in2 => \N__26775\,
            in3 => \N__26844\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41176\,
            in1 => \N__26835\,
            in2 => \_gnd_net_\,
            in3 => \N__26807\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__27018\,
            sr => \N__47037\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28488\,
            in1 => \N__28452\,
            in2 => \_gnd_net_\,
            in3 => \N__41178\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__27018\,
            sr => \N__47037\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41177\,
            in1 => \N__40755\,
            in2 => \_gnd_net_\,
            in3 => \N__41242\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47454\,
            ce => \N__27018\,
            sr => \N__47037\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__31296\,
            in1 => \N__31319\,
            in2 => \N__27033\,
            in3 => \N__26694\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26693\,
            in1 => \N__31295\,
            in2 => \N__31323\,
            in3 => \N__27029\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26762\,
            in1 => \N__26718\,
            in2 => \_gnd_net_\,
            in3 => \N__41174\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47444\,
            ce => \N__27016\,
            sr => \N__47044\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41171\,
            in1 => \N__26662\,
            in2 => \_gnd_net_\,
            in3 => \N__26678\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => \elapsed_time_ns_1_RNIV0CN9_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__26663\,
            in1 => \_gnd_net_\,
            in2 => \N__26628\,
            in3 => \N__41173\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47444\,
            ce => \N__27016\,
            sr => \N__47044\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__41172\,
            in1 => \N__27102\,
            in2 => \_gnd_net_\,
            in3 => \N__27078\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47444\,
            ce => \N__27016\,
            sr => \N__47044\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__26994\,
            in1 => \N__31241\,
            in2 => \N__31274\,
            in3 => \N__26978\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__26967\,
            in1 => \N__28141\,
            in2 => \_gnd_net_\,
            in3 => \N__29733\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47439\,
            ce => 'H',
            sr => \N__47049\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40605\,
            in1 => \N__42755\,
            in2 => \N__40129\,
            in3 => \N__37134\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31638\,
            in1 => \N__29286\,
            in2 => \_gnd_net_\,
            in3 => \N__35276\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__35277\,
            in1 => \N__31626\,
            in2 => \_gnd_net_\,
            in3 => \N__29478\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31614\,
            in1 => \N__29469\,
            in2 => \_gnd_net_\,
            in3 => \N__35278\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26913\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47420\,
            ce => 'H',
            sr => \N__47082\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__27915\,
            in1 => \N__27494\,
            in2 => \_gnd_net_\,
            in3 => \N__35884\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__27495\,
            in1 => \N__27477\,
            in2 => \N__35902\,
            in3 => \N__27914\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_10_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__27459\,
            in1 => \N__27447\,
            in2 => \N__29881\,
            in3 => \N__27435\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_10_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__29868\,
            in1 => \N__27411\,
            in2 => \N__27399\,
            in3 => \N__27372\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_10_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001110010"
        )
    port map (
            in0 => \N__29867\,
            in1 => \N__27360\,
            in2 => \N__27348\,
            in3 => \N__27333\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__27309\,
            in1 => \N__27285\,
            in2 => \N__29880\,
            in3 => \N__27273\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_10_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__29866\,
            in1 => \N__27249\,
            in2 => \N__27237\,
            in3 => \N__27210\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_10_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27198\,
            in2 => \N__27180\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_10_26_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_10_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27153\,
            in2 => \N__27135\,
            in3 => \N__27105\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_10_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27831\,
            in2 => \N__27813\,
            in3 => \N__27792\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_10_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27789\,
            in2 => \N__27774\,
            in3 => \N__27741\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27738\,
            in2 => \N__27720\,
            in3 => \N__27693\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_10_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27690\,
            in2 => \N__27672\,
            in3 => \N__27645\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27642\,
            in2 => \N__27624\,
            in3 => \N__27600\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_10_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27597\,
            in2 => \N__27585\,
            in3 => \N__27561\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_10_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27558\,
            in2 => \N__27543\,
            in3 => \N__27516\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_10_27_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_10_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27513\,
            in2 => \N__28095\,
            in3 => \N__28065\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_10_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27908\,
            in2 => \N__28062\,
            in3 => \N__28035\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27911\,
            in2 => \N__28032\,
            in3 => \N__28008\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_10_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27909\,
            in2 => \N__28005\,
            in3 => \N__27978\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27912\,
            in2 => \N__27975\,
            in3 => \N__27948\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27910\,
            in2 => \N__27945\,
            in3 => \N__27918\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27913\,
            in2 => \N__27870\,
            in3 => \N__27852\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27849\,
            in1 => \N__27843\,
            in2 => \_gnd_net_\,
            in3 => \N__27834\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29714\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29693\,
            ce => 'H',
            sr => \N__46975\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31830\,
            in2 => \N__29598\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32025\,
            in1 => \N__30071\,
            in2 => \_gnd_net_\,
            in3 => \N__28116\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32082\,
            in1 => \N__30159\,
            in2 => \N__30035\,
            in3 => \N__28113\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32026\,
            in1 => \N__29993\,
            in2 => \_gnd_net_\,
            in3 => \N__28110\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32083\,
            in1 => \N__29969\,
            in2 => \_gnd_net_\,
            in3 => \N__28107\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32027\,
            in1 => \N__30428\,
            in2 => \_gnd_net_\,
            in3 => \N__28104\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32084\,
            in1 => \N__30380\,
            in2 => \_gnd_net_\,
            in3 => \N__28101\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32028\,
            in1 => \N__30356\,
            in2 => \_gnd_net_\,
            in3 => \N__28098\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__47522\,
            ce => 'H',
            sr => \N__46981\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32017\,
            in1 => \N__30296\,
            in2 => \_gnd_net_\,
            in3 => \N__28209\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31956\,
            in1 => \N__30260\,
            in2 => \_gnd_net_\,
            in3 => \N__28206\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32014\,
            in1 => \N__30221\,
            in2 => \_gnd_net_\,
            in3 => \N__28203\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31957\,
            in1 => \N__30185\,
            in2 => \_gnd_net_\,
            in3 => \N__28200\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32015\,
            in1 => \N__30665\,
            in2 => \_gnd_net_\,
            in3 => \N__28197\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31958\,
            in1 => \N__30620\,
            in2 => \_gnd_net_\,
            in3 => \N__28194\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32016\,
            in1 => \N__30578\,
            in2 => \_gnd_net_\,
            in3 => \N__28191\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31959\,
            in1 => \N__28186\,
            in2 => \_gnd_net_\,
            in3 => \N__28170\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__47511\,
            ce => 'H',
            sr => \N__46989\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31960\,
            in1 => \N__28166\,
            in2 => \_gnd_net_\,
            in3 => \N__28149\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31964\,
            in1 => \N__28429\,
            in2 => \_gnd_net_\,
            in3 => \N__28413\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31961\,
            in1 => \N__28405\,
            in2 => \_gnd_net_\,
            in3 => \N__28389\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31965\,
            in1 => \N__28372\,
            in2 => \_gnd_net_\,
            in3 => \N__28356\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31962\,
            in1 => \N__28348\,
            in2 => \_gnd_net_\,
            in3 => \N__28326\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31966\,
            in1 => \N__28318\,
            in2 => \_gnd_net_\,
            in3 => \N__28302\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31963\,
            in1 => \N__28294\,
            in2 => \_gnd_net_\,
            in3 => \N__28275\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31967\,
            in1 => \N__28270\,
            in2 => \_gnd_net_\,
            in3 => \N__28254\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__47497\,
            ce => 'H',
            sr => \N__46998\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32050\,
            in1 => \N__28246\,
            in2 => \_gnd_net_\,
            in3 => \N__28230\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32067\,
            in1 => \N__28225\,
            in2 => \_gnd_net_\,
            in3 => \N__28566\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32051\,
            in1 => \N__28555\,
            in2 => \_gnd_net_\,
            in3 => \N__28536\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32068\,
            in1 => \N__28533\,
            in2 => \_gnd_net_\,
            in3 => \N__28518\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32052\,
            in1 => \N__28514\,
            in2 => \_gnd_net_\,
            in3 => \N__28497\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32069\,
            in1 => \N__28677\,
            in2 => \_gnd_net_\,
            in3 => \N__28494\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32053\,
            in1 => \N__28646\,
            in2 => \_gnd_net_\,
            in3 => \N__28491\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47485\,
            ce => 'H',
            sr => \N__47006\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28486\,
            in1 => \N__28445\,
            in2 => \_gnd_net_\,
            in3 => \N__40952\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011010100"
        )
    port map (
            in0 => \N__28658\,
            in1 => \N__28641\,
            in2 => \N__28625\,
            in3 => \N__28674\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28487\,
            in1 => \N__28444\,
            in2 => \_gnd_net_\,
            in3 => \N__40954\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47472\,
            ce => \N__32081\,
            sr => \N__47011\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011011101"
        )
    port map (
            in0 => \N__28659\,
            in1 => \N__28645\,
            in2 => \N__28626\,
            in3 => \N__28676\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__40953\,
            in1 => \N__40751\,
            in2 => \_gnd_net_\,
            in3 => \N__41243\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47472\,
            ce => \N__32081\,
            sr => \N__47011\
        );

    \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__28675\,
            in1 => \N__28657\,
            in2 => \N__28647\,
            in3 => \N__28621\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__30136\,
            in1 => \N__30782\,
            in2 => \N__28608\,
            in3 => \N__30771\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011111101"
        )
    port map (
            in0 => \N__31494\,
            in1 => \N__28605\,
            in2 => \N__31467\,
            in3 => \N__28589\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32275\,
            in2 => \_gnd_net_\,
            in3 => \N__28799\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__31492\,
            in1 => \N__28603\,
            in2 => \N__31466\,
            in3 => \N__28585\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__28604\,
            in1 => \N__31462\,
            in2 => \N__28590\,
            in3 => \N__31493\,
            lcout => OPEN,
            ltout => \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__32228\,
            in1 => \N__29162\,
            in2 => \N__28572\,
            in3 => \N__29151\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28569\,
            in3 => \N__32274\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__32276\,
            in1 => \N__32470\,
            in2 => \N__28803\,
            in3 => \N__30740\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47462\,
            ce => 'H',
            sr => \N__47018\
        );

    \phase_controller_inst2.stoper_hc.running_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__32229\,
            in1 => \N__32249\,
            in2 => \N__32315\,
            in3 => \N__32277\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47462\,
            ce => 'H',
            sr => \N__47018\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28791\,
            in2 => \N__28779\,
            in3 => \N__30736\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28770\,
            in2 => \N__28764\,
            in3 => \N__30719\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30695\,
            in1 => \N__28755\,
            in2 => \N__28746\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30680\,
            in1 => \N__28734\,
            in2 => \N__28725\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28716\,
            in2 => \N__28710\,
            in3 => \N__30965\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28698\,
            in2 => \N__28686\,
            in3 => \N__30950\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30935\,
            in1 => \N__28947\,
            in2 => \N__28938\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28929\,
            in2 => \N__28917\,
            in3 => \N__30920\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28908\,
            in2 => \N__28902\,
            in3 => \N__30905\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28893\,
            in2 => \N__28881\,
            in3 => \N__30890\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28872\,
            in2 => \N__28866\,
            in3 => \N__30875\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28857\,
            in2 => \N__28851\,
            in3 => \N__30860\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28830\,
            in2 => \N__28842\,
            in3 => \N__31160\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28821\,
            in2 => \N__28812\,
            in3 => \N__31145\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31130\,
            in1 => \N__29100\,
            in2 => \N__29112\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29094\,
            in2 => \N__29082\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29067\,
            in2 => \N__29055\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29040\,
            in2 => \N__29031\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29019\,
            in2 => \N__29010\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28995\,
            in2 => \N__28989\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28977\,
            in2 => \N__28971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28962\,
            in2 => \N__28956\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29181\,
            in2 => \N__29169\,
            in3 => \N__29142\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29139\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29136\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31755\,
            in2 => \_gnd_net_\,
            in3 => \N__31432\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29121\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47434\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__29202\,
            in1 => \N__33151\,
            in2 => \N__33468\,
            in3 => \N__32699\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47430\,
            ce => 'H',
            sr => \N__47050\
        );

    \phase_controller_inst1.state_3_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__31760\,
            in1 => \N__46388\,
            in2 => \N__31437\,
            in3 => \N__35786\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47430\,
            ce => 'H',
            sr => \N__47050\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__40128\,
            in1 => \N__40585\,
            in2 => \N__42852\,
            in3 => \N__37164\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__43139\,
            in1 => \N__40126\,
            in2 => \N__40626\,
            in3 => \N__37379\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \N__40125\,
            in1 => \N__37067\,
            in2 => \N__42672\,
            in3 => \N__40587\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40583\,
            in1 => \N__40121\,
            in2 => \N__46275\,
            in3 => \N__36885\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46373\,
            in1 => \N__40586\,
            in2 => \N__40229\,
            in3 => \N__37430\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40584\,
            in1 => \N__40127\,
            in2 => \N__42408\,
            in3 => \N__37547\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32700\,
            in2 => \_gnd_net_\,
            in3 => \N__29201\,
            lcout => \phase_controller_inst1.state_RNI7NN7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000101"
        )
    port map (
            in0 => \N__43281\,
            in1 => \N__38315\,
            in2 => \N__40627\,
            in3 => \N__40120\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32925\,
            in2 => \N__33057\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32797\,
            in2 => \N__31386\,
            in3 => \N__39444\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39445\,
            in1 => \N__39785\,
            in2 => \N__29190\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39800\,
            in2 => \N__31416\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39786\,
            in2 => \N__31395\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39801\,
            in2 => \N__29241\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39787\,
            in2 => \N__31512\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39802\,
            in2 => \N__29229\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39819\,
            in2 => \N__34632\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29217\,
            in2 => \N__39972\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39823\,
            in2 => \N__34728\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29211\,
            in2 => \N__39973\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39827\,
            in2 => \N__29277\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31404\,
            in2 => \N__39974\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39831\,
            in2 => \N__34602\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29265\,
            in2 => \N__39975\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39976\,
            in2 => \N__34713\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34839\,
            in2 => \N__40133\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39980\,
            in2 => \N__34686\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34827\,
            in2 => \N__40134\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39984\,
            in2 => \N__37287\,
            in3 => \N__29244\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34815\,
            in2 => \N__40135\,
            in3 => \N__29355\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39988\,
            in2 => \N__39345\,
            in3 => \N__29340\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34698\,
            in2 => \N__40136\,
            in3 => \N__29325\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40008\,
            in2 => \N__34659\,
            in3 => \N__29322\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_11_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34803\,
            in2 => \N__40141\,
            in3 => \N__29307\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40012\,
            in2 => \N__37395\,
            in3 => \N__29304\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32943\,
            in2 => \N__40142\,
            in3 => \N__29289\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40016\,
            in2 => \N__34776\,
            in3 => \N__29280\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29487\,
            in2 => \N__40143\,
            in3 => \N__29472\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40020\,
            in2 => \N__39387\,
            in3 => \N__29463\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__32964\,
            in1 => \N__31599\,
            in2 => \N__35296\,
            in3 => \N__29460\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__35283\,
            in1 => \_gnd_net_\,
            in2 => \N__31665\,
            in3 => \N__29445\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__31533\,
            in1 => \N__29424\,
            in2 => \_gnd_net_\,
            in3 => \N__35282\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S1_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39603\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47417\,
            ce => 'H',
            sr => \N__47077\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_11_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29388\,
            in2 => \N__29886\,
            in3 => \N__29885\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_11_24_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_11_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29382\,
            in2 => \_gnd_net_\,
            in3 => \N__29370\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_11_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29895\,
            in2 => \_gnd_net_\,
            in3 => \N__29580\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29577\,
            in2 => \_gnd_net_\,
            in3 => \N__29571\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29568\,
            in2 => \_gnd_net_\,
            in3 => \N__29562\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_11_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29742\,
            in2 => \_gnd_net_\,
            in3 => \N__29559\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29556\,
            in2 => \_gnd_net_\,
            in3 => \N__29550\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_11_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29547\,
            in2 => \_gnd_net_\,
            in3 => \N__29541\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_11_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29538\,
            in2 => \_gnd_net_\,
            in3 => \N__29526\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_11_25_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_11_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__29523\,
            in1 => \N__29511\,
            in2 => \N__29872\,
            in3 => \N__29499\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_11_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111110000"
        )
    port map (
            in0 => \N__29496\,
            in1 => \N__29937\,
            in2 => \N__29916\,
            in3 => \N__29829\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__29830\,
            in1 => \N__29793\,
            in2 => \N__29784\,
            in3 => \N__29760\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29713\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29694\,
            ce => 'H',
            sr => \N__46969\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29682\,
            in1 => \N__29636\,
            in2 => \_gnd_net_\,
            in3 => \N__41168\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47509\,
            ce => \N__32029\,
            sr => \N__46976\
        );

    \phase_controller_inst1.start_timer_hc_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__46466\,
            in1 => \N__30153\,
            in2 => \N__33131\,
            in3 => \N__29613\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47496\,
            ce => 'H',
            sr => \N__46982\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47496\,
            ce => 'H',
            sr => \N__46982\
        );

    \phase_controller_inst1.stoper_hc.running_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111100001010"
        )
    port map (
            in0 => \N__32158\,
            in1 => \N__30758\,
            in2 => \N__30137\,
            in3 => \N__29589\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47496\,
            ce => 'H',
            sr => \N__46982\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32157\,
            in2 => \_gnd_net_\,
            in3 => \N__32137\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__30128\,
            in1 => \N__29588\,
            in2 => \_gnd_net_\,
            in3 => \N__30150\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30162\,
            in3 => \N__32138\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011100100"
        )
    port map (
            in0 => \N__32159\,
            in1 => \N__32731\,
            in2 => \N__30138\,
            in3 => \N__30759\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47496\,
            ce => 'H',
            sr => \N__46982\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__30151\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30129\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30105\,
            in2 => \N__30093\,
            in3 => \N__31822\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_12_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30084\,
            in2 => \N__30057\,
            in3 => \N__30072\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30048\,
            in2 => \N__30015\,
            in3 => \N__30036\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30006\,
            in2 => \N__29979\,
            in3 => \N__29994\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29970\,
            in1 => \N__29955\,
            in2 => \N__29946\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30429\,
            in1 => \N__30414\,
            in2 => \N__30402\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30390\,
            in2 => \N__30366\,
            in3 => \N__30381\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30357\,
            in1 => \N__30342\,
            in2 => \N__30324\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30312\,
            in2 => \N__30282\,
            in3 => \N__30300\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_12_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30273\,
            in2 => \N__30246\,
            in3 => \N__30261\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30237\,
            in2 => \N__30207\,
            in3 => \N__30225\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30195\,
            in2 => \N__30171\,
            in3 => \N__30186\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30666\,
            in1 => \N__30651\,
            in2 => \N__30636\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30624\,
            in1 => \N__30594\,
            in2 => \N__30606\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30588\,
            in2 => \N__30564\,
            in3 => \N__30579\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30555\,
            in2 => \N__30546\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30531\,
            in2 => \N__30519\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30504\,
            in2 => \N__30495\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30483\,
            in2 => \N__30471\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30456\,
            in2 => \N__30444\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30846\,
            in2 => \N__30834\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30819\,
            in2 => \N__30807\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30792\,
            in2 => \N__30786\,
            in3 => \N__30765\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30762\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30747\,
            in2 => \N__30741\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32455\,
            in1 => \N__30720\,
            in2 => \_gnd_net_\,
            in3 => \N__30708\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__32459\,
            in1 => \N__30696\,
            in2 => \N__30705\,
            in3 => \N__30684\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32456\,
            in1 => \N__30681\,
            in2 => \_gnd_net_\,
            in3 => \N__30669\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32460\,
            in1 => \N__30966\,
            in2 => \_gnd_net_\,
            in3 => \N__30954\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32457\,
            in1 => \N__30951\,
            in2 => \_gnd_net_\,
            in3 => \N__30939\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32461\,
            in1 => \N__30936\,
            in2 => \_gnd_net_\,
            in3 => \N__30924\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32458\,
            in1 => \N__30921\,
            in2 => \_gnd_net_\,
            in3 => \N__30909\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__47453\,
            ce => 'H',
            sr => \N__47012\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32450\,
            in1 => \N__30906\,
            in2 => \_gnd_net_\,
            in3 => \N__30894\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32462\,
            in1 => \N__30891\,
            in2 => \_gnd_net_\,
            in3 => \N__30879\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32447\,
            in1 => \N__30876\,
            in2 => \_gnd_net_\,
            in3 => \N__30864\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32463\,
            in1 => \N__30861\,
            in2 => \_gnd_net_\,
            in3 => \N__30849\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32448\,
            in1 => \N__31161\,
            in2 => \_gnd_net_\,
            in3 => \N__31149\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32464\,
            in1 => \N__31146\,
            in2 => \_gnd_net_\,
            in3 => \N__31134\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32449\,
            in1 => \N__31131\,
            in2 => \_gnd_net_\,
            in3 => \N__31119\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32465\,
            in1 => \N__31106\,
            in2 => \_gnd_net_\,
            in3 => \N__31092\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__47443\,
            ce => 'H',
            sr => \N__47019\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32451\,
            in1 => \N__31087\,
            in2 => \_gnd_net_\,
            in3 => \N__31071\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32466\,
            in1 => \N__31061\,
            in2 => \_gnd_net_\,
            in3 => \N__31047\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32452\,
            in1 => \N__31034\,
            in2 => \_gnd_net_\,
            in3 => \N__31020\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32467\,
            in1 => \N__31010\,
            in2 => \_gnd_net_\,
            in3 => \N__30996\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32453\,
            in1 => \N__30983\,
            in2 => \_gnd_net_\,
            in3 => \N__30969\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32468\,
            in1 => \N__31364\,
            in2 => \_gnd_net_\,
            in3 => \N__31350\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32454\,
            in1 => \N__31340\,
            in2 => \_gnd_net_\,
            in3 => \N__31326\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32469\,
            in1 => \N__31313\,
            in2 => \_gnd_net_\,
            in3 => \N__31299\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__47438\,
            ce => 'H',
            sr => \N__47026\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32474\,
            in1 => \N__31294\,
            in2 => \_gnd_net_\,
            in3 => \N__31278\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32478\,
            in1 => \N__31267\,
            in2 => \_gnd_net_\,
            in3 => \N__31248\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32475\,
            in1 => \N__31237\,
            in2 => \_gnd_net_\,
            in3 => \N__31215\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32479\,
            in1 => \N__31202\,
            in2 => \_gnd_net_\,
            in3 => \N__31188\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32476\,
            in1 => \N__31178\,
            in2 => \_gnd_net_\,
            in3 => \N__31164\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32480\,
            in1 => \N__31491\,
            in2 => \_gnd_net_\,
            in3 => \N__31473\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32477\,
            in1 => \N__31451\,
            in2 => \_gnd_net_\,
            in3 => \N__31470\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47433\,
            ce => 'H',
            sr => \N__47032\
        );

    \phase_controller_inst1.state_2_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111000001010"
        )
    port map (
            in0 => \N__32714\,
            in1 => \N__31759\,
            in2 => \N__32754\,
            in3 => \N__31436\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47429\,
            ce => 'H',
            sr => \N__47038\
        );

    \phase_controller_inst1.state_RNIE87F_2_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32713\,
            in2 => \_gnd_net_\,
            in3 => \N__32749\,
            lcout => \phase_controller_inst1.state_RNIE87FZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40580\,
            in1 => \N__42487\,
            in2 => \N__40230\,
            in3 => \N__36848\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__39954\,
            in1 => \N__40576\,
            in2 => \N__37034\,
            in3 => \N__42621\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40573\,
            in1 => \N__39956\,
            in2 => \N__42453\,
            in3 => \N__36816\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__37472\,
            in1 => \N__40571\,
            in2 => \N__32807\,
            in3 => \N__39498\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40575\,
            in1 => \N__39958\,
            in2 => \N__42851\,
            in3 => \N__37163\,
            lcout => \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__39955\,
            in1 => \N__40572\,
            in2 => \N__42495\,
            in3 => \N__36849\,
            lcout => \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40574\,
            in1 => \N__39957\,
            in2 => \N__42360\,
            in3 => \N__37196\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32921\,
            in2 => \N__32892\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32796\,
            in2 => \N__32775\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32625\,
            in2 => \N__39965\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39791\,
            in2 => \N__31503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32847\,
            in2 => \N__39966\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39795\,
            in2 => \N__32841\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32832\,
            in2 => \N__39967\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39799\,
            in2 => \N__31524\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39803\,
            in2 => \N__32826\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32910\,
            in2 => \N__39968\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39807\,
            in2 => \N__32817\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32982\,
            in2 => \N__39969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39811\,
            in2 => \N__32871\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32904\,
            in2 => \N__39970\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39815\,
            in2 => \N__34617\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32862\,
            in2 => \N__39971\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32898\,
            in2 => \N__40137\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39995\,
            in2 => \N__32856\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32877\,
            in2 => \N__40138\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39999\,
            in2 => \N__34791\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34671\,
            in2 => \N__40139\,
            in3 => \N__31581\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40003\,
            in2 => \N__32952\,
            in3 => \N__31566\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38088\,
            in2 => \N__40140\,
            in3 => \N__31551\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40007\,
            in2 => \N__37272\,
            in3 => \N__31536\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40021\,
            in2 => \N__37323\,
            in3 => \N__31527\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37809\,
            in2 => \N__40144\,
            in3 => \N__31668\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40025\,
            in2 => \N__39663\,
            in3 => \N__31656\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32934\,
            in2 => \N__40145\,
            in3 => \N__31641\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40029\,
            in2 => \N__32976\,
            in3 => \N__31629\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38289\,
            in2 => \N__40146\,
            in3 => \N__31617\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40033\,
            in2 => \N__37338\,
            in3 => \N__31605\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__40034\,
            in1 => \N__40444\,
            in2 => \_gnd_net_\,
            in3 => \N__31602\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.stop_timer_s1_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__31784\,
            in1 => \N__31769\,
            in2 => \N__33024\,
            in3 => \N__33041\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47419\,
            ce => 'H',
            sr => \N__47065\
        );

    \current_shift_inst.timer_s1.running_LC_12_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__33042\,
            in1 => \N__33020\,
            in2 => \_gnd_net_\,
            in3 => \N__41306\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47419\,
            ce => 'H',
            sr => \N__47065\
        );

    \phase_controller_inst1.S1_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31770\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47419\,
            ce => 'H',
            sr => \N__47065\
        );

    \current_shift_inst.start_timer_s1_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__31783\,
            in1 => \N__33040\,
            in2 => \_gnd_net_\,
            in3 => \N__31768\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47419\,
            ce => 'H',
            sr => \N__47065\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_12_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__35839\,
            in1 => \N__36078\,
            in2 => \N__36000\,
            in3 => \N__31734\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__36079\,
            in1 => \N__35840\,
            in2 => \N__31728\,
            in3 => \N__35950\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_12_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010011"
        )
    port map (
            in0 => \N__35841\,
            in1 => \N__36080\,
            in2 => \N__36001\,
            in3 => \N__31719\,
            lcout => \pwm_generator_inst.un14_counter_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_12_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__36081\,
            in1 => \N__35951\,
            in2 => \N__31713\,
            in3 => \N__35842\,
            lcout => \pwm_generator_inst.un14_counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_12_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__36075\,
            in1 => \N__35939\,
            in2 => \N__31704\,
            in3 => \N__35836\,
            lcout => \pwm_generator_inst.un14_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__35838\,
            in1 => \N__36077\,
            in2 => \N__35999\,
            in3 => \N__31695\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_12_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__36076\,
            in1 => \N__35943\,
            in2 => \N__31689\,
            in3 => \N__35837\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001111"
        )
    port map (
            in0 => \N__35852\,
            in1 => \N__32187\,
            in2 => \N__36090\,
            in3 => \N__35953\,
            lcout => \pwm_generator_inst.un14_counter_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_12_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__35952\,
            in1 => \N__35853\,
            in2 => \N__32181\,
            in3 => \N__36088\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__47121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pll_inst.red_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_1_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__35731\,
            in1 => \N__41927\,
            in2 => \_gnd_net_\,
            in3 => \N__35709\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47543\,
            ce => 'H',
            sr => \N__46959\
        );

    \phase_controller_inst2.start_timer_hc_RNO_0_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39576\,
            lcout => \phase_controller_inst2.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44706\,
            in1 => \N__44321\,
            in2 => \_gnd_net_\,
            in3 => \N__48332\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47523\,
            ce => \N__47825\,
            sr => \N__46970\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__46563\,
            in1 => \N__36945\,
            in2 => \N__38854\,
            in3 => \N__47874\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47512\,
            ce => 'H',
            sr => \N__46977\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__32160\,
            in1 => \N__31826\,
            in2 => \N__32142\,
            in3 => \N__31984\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47512\,
            ce => 'H',
            sr => \N__46977\
        );

    \phase_controller_inst2.start_timer_hc_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__31806\,
            in1 => \N__46456\,
            in2 => \N__32295\,
            in3 => \N__35708\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47512\,
            ce => 'H',
            sr => \N__46977\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32215\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32290\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32294\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47512\,
            ce => 'H',
            sr => \N__46977\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__32214\,
            in1 => \N__32319\,
            in2 => \_gnd_net_\,
            in3 => \N__32289\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst2.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000001010"
        )
    port map (
            in0 => \N__38122\,
            in1 => \N__32256\,
            in2 => \N__32232\,
            in3 => \N__32216\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47512\,
            ce => 'H',
            sr => \N__46977\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33380\,
            in2 => \N__36231\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33353\,
            in2 => \N__33414\,
            in3 => \N__32199\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33332\,
            in2 => \N__33384\,
            in3 => \N__32196\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33354\,
            in2 => \N__33719\,
            in3 => \N__32193\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33333\,
            in2 => \N__33692\,
            in3 => \N__32190\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33659\,
            in2 => \N__33720\,
            in3 => \N__32514\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33625\,
            in2 => \N__33693\,
            in3 => \N__32511\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33595\,
            in2 => \N__33663\,
            in3 => \N__32508\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__47498\,
            ce => \N__36196\,
            sr => \N__46983\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33633\,
            in2 => \N__33575\,
            in3 => \N__32505\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33548\,
            in2 => \N__33606\,
            in3 => \N__32502\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33527\,
            in2 => \N__33576\,
            in3 => \N__32499\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33549\,
            in2 => \N__33938\,
            in3 => \N__32496\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33528\,
            in2 => \N__33911\,
            in3 => \N__32493\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33881\,
            in2 => \N__33939\,
            in3 => \N__32490\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33844\,
            in2 => \N__33912\,
            in3 => \N__32541\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33814\,
            in2 => \N__33882\,
            in3 => \N__32538\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__47486\,
            ce => \N__36195\,
            sr => \N__46990\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33794\,
            in2 => \N__33852\,
            in3 => \N__32535\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33770\,
            in2 => \N__33825\,
            in3 => \N__32532\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33795\,
            in2 => \N__33749\,
            in3 => \N__32529\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33771\,
            in2 => \N__34217\,
            in3 => \N__32526\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34190\,
            in2 => \N__33750\,
            in3 => \N__32523\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34169\,
            in2 => \N__34218\,
            in3 => \N__32520\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34191\,
            in2 => \N__34139\,
            in3 => \N__32517\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34099\,
            in2 => \N__34170\,
            in3 => \N__32562\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__47473\,
            ce => \N__36194\,
            sr => \N__46999\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34140\,
            in2 => \N__34079\,
            in3 => \N__32559\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__47463\,
            ce => \N__36178\,
            sr => \N__47007\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34052\,
            in2 => \N__34110\,
            in3 => \N__32556\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__47463\,
            ce => \N__36178\,
            sr => \N__47007\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34032\,
            in2 => \N__34080\,
            in3 => \N__32553\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__47463\,
            ce => \N__36178\,
            sr => \N__47007\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34053\,
            in2 => \N__34011\,
            in3 => \N__32550\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__47463\,
            ce => \N__36178\,
            sr => \N__47007\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32547\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47463\,
            ce => \N__36178\,
            sr => \N__47007\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__39066\,
            in1 => \N__39089\,
            in2 => \N__32619\,
            in3 => \N__32604\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__32603\,
            in1 => \N__39065\,
            in2 => \N__39093\,
            in3 => \N__32615\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36292\,
            in1 => \N__36305\,
            in2 => \_gnd_net_\,
            in3 => \N__48263\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => \elapsed_time_ns_1_RNI1CPBB_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__48266\,
            in1 => \N__36293\,
            in2 => \N__32544\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47455\,
            ce => \N__47875\,
            sr => \N__47013\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36369\,
            in1 => \N__48264\,
            in2 => \_gnd_net_\,
            in3 => \N__36332\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48265\,
            in1 => \_gnd_net_\,
            in2 => \N__32607\,
            in3 => \N__36370\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47455\,
            ce => \N__47875\,
            sr => \N__47013\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45340\,
            in1 => \N__45378\,
            in2 => \_gnd_net_\,
            in3 => \N__48267\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47455\,
            ce => \N__47875\,
            sr => \N__47013\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__32590\,
            in1 => \N__39232\,
            in2 => \N__39272\,
            in3 => \N__32578\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48333\,
            in1 => \N__41833\,
            in2 => \_gnd_net_\,
            in3 => \N__41798\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => \elapsed_time_ns_1_RNIVAQBB_0_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__41834\,
            in1 => \_gnd_net_\,
            in2 => \N__32595\,
            in3 => \N__48335\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47445\,
            ce => \N__47877\,
            sr => \N__47020\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__32580\,
            in1 => \N__32592\,
            in2 => \N__39237\,
            in3 => \N__39271\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__32591\,
            in1 => \N__39233\,
            in2 => \N__39273\,
            in3 => \N__32579\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48334\,
            in1 => \N__46172\,
            in2 => \_gnd_net_\,
            in3 => \N__46146\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47445\,
            ce => \N__47877\,
            sr => \N__47020\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33078\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43170\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__43229\,
            sr => \N__47027\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47440\,
            ce => \N__43229\,
            sr => \N__47027\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38005\,
            in1 => \N__36912\,
            in2 => \_gnd_net_\,
            in3 => \N__33079\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42576\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__33155\,
            in1 => \N__33461\,
            in2 => \N__32753\,
            in3 => \N__32715\,
            lcout => \phase_controller_inst1.start_timer_tr_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_ns_i_a3_1_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46433\,
            lcout => state_ns_i_a3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000011001100"
        )
    port map (
            in0 => \N__47576\,
            in1 => \N__32689\,
            in2 => \N__46656\,
            in3 => \N__46546\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47431\,
            ce => 'H',
            sr => \N__47039\
        );

    \phase_controller_inst1.state_4_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__46434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32653\,
            lcout => phase_controller_inst1_state_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47431\,
            ce => 'H',
            sr => \N__47039\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40577\,
            in1 => \N__46271\,
            in2 => \N__40231\,
            in3 => \N__36881\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__36815\,
            in1 => \N__40578\,
            in2 => \N__40232\,
            in3 => \N__42449\,
            lcout => \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38006\,
            in1 => \N__42488\,
            in2 => \_gnd_net_\,
            in3 => \N__36847\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__42399\,
            in1 => \N__40150\,
            in2 => \N__37548\,
            in3 => \N__40579\,
            lcout => \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40483\,
            in1 => \N__40112\,
            in2 => \N__42359\,
            in3 => \N__37197\,
            lcout => \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40113\,
            in1 => \N__40484\,
            in2 => \N__37584\,
            in3 => \N__42800\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__40486\,
            in1 => \N__37104\,
            in2 => \N__42714\,
            in3 => \N__40111\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38016\,
            in1 => \N__42445\,
            in2 => \_gnd_net_\,
            in3 => \N__36814\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__40482\,
            in1 => \N__37473\,
            in2 => \N__32808\,
            in3 => \N__39497\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__35507\,
            in1 => \N__32766\,
            in2 => \_gnd_net_\,
            in3 => \N__34757\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__32891\,
            in1 => \_gnd_net_\,
            in2 => \N__32928\,
            in3 => \N__35508\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__40114\,
            in1 => \N__40485\,
            in2 => \N__42756\,
            in3 => \N__37130\,
            lcout => \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__40448\,
            in1 => \N__40200\,
            in2 => \N__37038\,
            in3 => \N__42620\,
            lcout => \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40202\,
            in1 => \N__40450\,
            in2 => \N__37782\,
            in3 => \N__43088\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__40445\,
            in1 => \N__33096\,
            in2 => \_gnd_net_\,
            in3 => \N__33087\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40204\,
            in1 => \N__40452\,
            in2 => \N__37623\,
            in3 => \N__43007\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__40447\,
            in1 => \N__40199\,
            in2 => \N__37074\,
            in3 => \N__42671\,
            lcout => \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__40201\,
            in1 => \N__40449\,
            in2 => \N__43140\,
            in3 => \N__37380\,
            lcout => \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40451\,
            in1 => \N__40203\,
            in2 => \N__43050\,
            in3 => \N__37716\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__40198\,
            in1 => \N__40446\,
            in2 => \N__46377\,
            in3 => \N__37434\,
            lcout => \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40196\,
            in1 => \N__40442\,
            in2 => \N__37881\,
            in3 => \N__43320\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__40195\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40443\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40197\,
            in1 => \N__40441\,
            in2 => \N__37239\,
            in3 => \N__42893\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__37957\,
            in1 => \N__42892\,
            in2 => \_gnd_net_\,
            in3 => \N__37235\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47425\,
            ce => \N__43227\,
            sr => \N__47058\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40362\,
            in1 => \N__43352\,
            in2 => \N__40256\,
            in3 => \N__38072\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__43353\,
            in1 => \N__40363\,
            in2 => \N__38073\,
            in3 => \N__40208\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43193\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47422\,
            ce => \N__43226\,
            sr => \N__47061\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36924\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__33086\,
            in1 => \N__40361\,
            in2 => \N__33060\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__41302\,
            in1 => \N__33019\,
            in2 => \_gnd_net_\,
            in3 => \N__33039\,
            lcout => \current_shift_inst.timer_s1.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41301\,
            in2 => \_gnd_net_\,
            in3 => \N__33018\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35208\,
            in2 => \_gnd_net_\,
            in3 => \N__38276\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__35209\,
            in1 => \_gnd_net_\,
            in2 => \N__38280\,
            in3 => \N__38255\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_201_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34962\,
            in1 => \N__35102\,
            in2 => \_gnd_net_\,
            in3 => \N__32991\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_22_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_1_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34956\,
            in1 => \N__35036\,
            in2 => \_gnd_net_\,
            in3 => \N__32988\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_2_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34963\,
            in1 => \N__35123\,
            in2 => \_gnd_net_\,
            in3 => \N__32985\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_3_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34957\,
            in1 => \N__35060\,
            in2 => \_gnd_net_\,
            in3 => \N__33180\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_4_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34964\,
            in1 => \N__35081\,
            in2 => \_gnd_net_\,
            in3 => \N__33177\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_5_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34958\,
            in1 => \N__34984\,
            in2 => \_gnd_net_\,
            in3 => \N__33174\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_6_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34965\,
            in1 => \N__35008\,
            in2 => \_gnd_net_\,
            in3 => \N__33171\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_7_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34959\,
            in1 => \N__35144\,
            in2 => \_gnd_net_\,
            in3 => \N__33168\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__47421\,
            ce => 'H',
            sr => \N__47066\
        );

    \pwm_generator_inst.counter_8_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34961\,
            in1 => \N__35165\,
            in2 => \_gnd_net_\,
            in3 => \N__33165\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__47418\,
            ce => 'H',
            sr => \N__47070\
        );

    \pwm_generator_inst.counter_9_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35186\,
            in1 => \N__34960\,
            in2 => \_gnd_net_\,
            in3 => \N__33162\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47418\,
            ce => 'H',
            sr => \N__47070\
        );

    \phase_controller_inst1.state_1_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__33159\,
            in1 => \N__33453\,
            in2 => \_gnd_net_\,
            in3 => \N__33132\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47418\,
            ce => 'H',
            sr => \N__47070\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33102\,
            in2 => \N__35802\,
            in3 => \N__35103\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_13_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_13_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35037\,
            in1 => \N__33303\,
            in2 => \N__33312\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33285\,
            in2 => \N__33297\,
            in3 => \N__35124\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33267\,
            in2 => \N__33279\,
            in3 => \N__35061\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35082\,
            in1 => \N__33249\,
            in2 => \N__33261\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33234\,
            in2 => \N__33243\,
            in3 => \N__34986\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_13_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35010\,
            in1 => \N__33219\,
            in2 => \N__33228\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_13_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33204\,
            in2 => \N__33213\,
            in3 => \N__35145\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33186\,
            in2 => \N__33198\,
            in3 => \N__35166\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_13_25_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33498\,
            in2 => \N__33507\,
            in3 => \N__35187\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_13_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33492\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47416\,
            ce => 'H',
            sr => \N__47078\
        );

    \phase_controller_inst1.S2_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33457\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47412\,
            ce => 'H',
            sr => \N__47092\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33407\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47544\,
            ce => \N__36204\,
            sr => \N__46960\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34343\,
            in1 => \N__36220\,
            in2 => \_gnd_net_\,
            in3 => \N__33417\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34347\,
            in1 => \N__33406\,
            in2 => \_gnd_net_\,
            in3 => \N__33387\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34344\,
            in1 => \N__33379\,
            in2 => \_gnd_net_\,
            in3 => \N__33357\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34348\,
            in1 => \N__33352\,
            in2 => \_gnd_net_\,
            in3 => \N__33336\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34345\,
            in1 => \N__33331\,
            in2 => \_gnd_net_\,
            in3 => \N__33315\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34349\,
            in1 => \N__33712\,
            in2 => \_gnd_net_\,
            in3 => \N__33696\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34346\,
            in1 => \N__33680\,
            in2 => \_gnd_net_\,
            in3 => \N__33666\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34350\,
            in1 => \N__33652\,
            in2 => \_gnd_net_\,
            in3 => \N__33636\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__47533\,
            ce => \N__33993\,
            sr => \N__46964\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34342\,
            in1 => \N__33626\,
            in2 => \_gnd_net_\,
            in3 => \N__33609\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34338\,
            in1 => \N__33599\,
            in2 => \_gnd_net_\,
            in3 => \N__33579\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34339\,
            in1 => \N__33568\,
            in2 => \_gnd_net_\,
            in3 => \N__33552\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34335\,
            in1 => \N__33547\,
            in2 => \_gnd_net_\,
            in3 => \N__33531\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34340\,
            in1 => \N__33526\,
            in2 => \_gnd_net_\,
            in3 => \N__33510\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34336\,
            in1 => \N__33931\,
            in2 => \_gnd_net_\,
            in3 => \N__33915\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34341\,
            in1 => \N__33899\,
            in2 => \_gnd_net_\,
            in3 => \N__33885\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34337\,
            in1 => \N__33874\,
            in2 => \_gnd_net_\,
            in3 => \N__33855\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__47524\,
            ce => \N__33992\,
            sr => \N__46971\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34307\,
            in1 => \N__33845\,
            in2 => \_gnd_net_\,
            in3 => \N__33828\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34331\,
            in1 => \N__33818\,
            in2 => \_gnd_net_\,
            in3 => \N__33798\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34308\,
            in1 => \N__33793\,
            in2 => \_gnd_net_\,
            in3 => \N__33774\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34332\,
            in1 => \N__33769\,
            in2 => \_gnd_net_\,
            in3 => \N__33753\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34309\,
            in1 => \N__33737\,
            in2 => \_gnd_net_\,
            in3 => \N__33723\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34333\,
            in1 => \N__34210\,
            in2 => \_gnd_net_\,
            in3 => \N__34194\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34310\,
            in1 => \N__34189\,
            in2 => \_gnd_net_\,
            in3 => \N__34173\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34334\,
            in1 => \N__34162\,
            in2 => \_gnd_net_\,
            in3 => \N__34143\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__47513\,
            ce => \N__33991\,
            sr => \N__46978\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34303\,
            in1 => \N__34135\,
            in2 => \_gnd_net_\,
            in3 => \N__34113\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__47499\,
            ce => \N__33984\,
            sr => \N__46984\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34311\,
            in1 => \N__34103\,
            in2 => \_gnd_net_\,
            in3 => \N__34083\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__47499\,
            ce => \N__33984\,
            sr => \N__46984\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34304\,
            in1 => \N__34072\,
            in2 => \_gnd_net_\,
            in3 => \N__34056\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__47499\,
            ce => \N__33984\,
            sr => \N__46984\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34312\,
            in1 => \N__34051\,
            in2 => \_gnd_net_\,
            in3 => \N__34035\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__47499\,
            ce => \N__33984\,
            sr => \N__46984\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__34305\,
            in1 => \N__34031\,
            in2 => \_gnd_net_\,
            in3 => \N__34017\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__47499\,
            ce => \N__33984\,
            sr => \N__46984\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34007\,
            in1 => \N__34306\,
            in2 => \_gnd_net_\,
            in3 => \N__34014\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47499\,
            ce => \N__33984\,
            sr => \N__46984\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35214\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48288\,
            in1 => \N__48426\,
            in2 => \_gnd_net_\,
            in3 => \N__48463\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47487\,
            ce => \N__47861\,
            sr => \N__46991\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45015\,
            in1 => \N__48291\,
            in2 => \_gnd_net_\,
            in3 => \N__44983\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47487\,
            ce => \N__47861\,
            sr => \N__46991\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44871\,
            in1 => \N__48292\,
            in2 => \_gnd_net_\,
            in3 => \N__36611\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47487\,
            ce => \N__47861\,
            sr => \N__46991\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48289\,
            in1 => \N__45084\,
            in2 => \_gnd_net_\,
            in3 => \N__45056\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47487\,
            ce => \N__47861\,
            sr => \N__46991\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44830\,
            in1 => \N__48290\,
            in2 => \_gnd_net_\,
            in3 => \N__36255\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47487\,
            ce => \N__47861\,
            sr => \N__46991\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__42277\,
            in1 => \N__41698\,
            in2 => \N__46147\,
            in3 => \N__36652\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34224\,
            in1 => \N__34401\,
            in2 => \N__34227\,
            in3 => \N__34407\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48358\,
            in1 => \N__45520\,
            in2 => \N__45767\,
            in3 => \N__41832\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36736\,
            in1 => \N__45301\,
            in2 => \N__44286\,
            in3 => \N__45181\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46487\,
            in1 => \N__36283\,
            in2 => \N__36375\,
            in3 => \N__45132\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__45133\,
            in1 => \N__48336\,
            in2 => \N__45116\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => \elapsed_time_ns_1_RNIV9PBB_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48337\,
            in1 => \_gnd_net_\,
            in2 => \N__34395\,
            in3 => \N__45134\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47474\,
            ce => \N__47876\,
            sr => \N__47000\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36495\,
            in2 => \N__34392\,
            in3 => \N__38855\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34383\,
            in2 => \N__36438\,
            in3 => \N__38823\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36381\,
            in2 => \N__34377\,
            in3 => \N__38793\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38772\,
            in1 => \N__44586\,
            in2 => \N__34368\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35688\,
            in2 => \N__34359\,
            in3 => \N__38754\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36243\,
            in2 => \N__34548\,
            in3 => \N__38736\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39042\,
            in1 => \N__34536\,
            in2 => \N__34527\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34518\,
            in2 => \N__34506\,
            in3 => \N__39024\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34497\,
            in2 => \N__34488\,
            in3 => \N__39006\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_14_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34467\,
            in2 => \N__34479\,
            in3 => \N__38988\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34461\,
            in2 => \N__34452\,
            in3 => \N__38970\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34440\,
            in2 => \N__34431\,
            in3 => \N__38952\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38934\,
            in1 => \N__34413\,
            in2 => \N__34422\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38916\,
            in1 => \N__36762\,
            in2 => \N__34587\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42252\,
            in2 => \N__34578\,
            in3 => \N__39210\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36708\,
            in2 => \N__36690\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42174\,
            in2 => \N__42318\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36549\,
            in2 => \N__36588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34569\,
            in2 => \N__34560\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45819\,
            in2 => \N__45882\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42162\,
            in2 => \N__45894\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46053\,
            in2 => \N__45990\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34644\,
            in2 => \N__36984\,
            in3 => \N__34638\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34635\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42345\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38002\,
            in1 => \N__46267\,
            in2 => \_gnd_net_\,
            in3 => \N__36868\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42838\,
            in1 => \N__38004\,
            in2 => \_gnd_net_\,
            in3 => \N__37151\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40598\,
            in1 => \N__40265\,
            in2 => \N__42801\,
            in3 => \N__37573\,
            lcout => \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40264\,
            in1 => \N__40600\,
            in2 => \N__37500\,
            in3 => \N__42577\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40599\,
            in1 => \N__40263\,
            in2 => \N__42582\,
            in3 => \N__37498\,
            lcout => \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42346\,
            in1 => \N__38003\,
            in2 => \_gnd_net_\,
            in3 => \N__37183\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__42710\,
            in1 => \N__40601\,
            in2 => \N__37100\,
            in3 => \N__40260\,
            lcout => \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38007\,
            in1 => \N__42709\,
            in2 => \_gnd_net_\,
            in3 => \N__37093\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__37774\,
            in1 => \N__40261\,
            in2 => \N__43095\,
            in3 => \N__40602\,
            lcout => \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40604\,
            in1 => \N__46319\,
            in2 => \N__40272\,
            in3 => \N__37681\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42670\,
            in1 => \N__38009\,
            in2 => \_gnd_net_\,
            in3 => \N__37054\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38010\,
            in1 => \N__42613\,
            in2 => \_gnd_net_\,
            in3 => \N__37015\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__37615\,
            in1 => \N__40262\,
            in2 => \N__43008\,
            in3 => \N__40603\,
            lcout => \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__38008\,
            in1 => \N__37118\,
            in2 => \_gnd_net_\,
            in3 => \N__42742\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42933\,
            in1 => \N__40615\,
            in2 => \N__40237\,
            in3 => \N__37654\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40617\,
            in1 => \N__43472\,
            in2 => \N__40234\,
            in3 => \N__37915\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43042\,
            in1 => \N__40612\,
            in2 => \N__40238\,
            in3 => \N__37708\,
            lcout => \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40613\,
            in1 => \N__42965\,
            in2 => \N__40235\,
            in3 => \N__37741\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__37234\,
            in1 => \N__42894\,
            in2 => \N__40236\,
            in3 => \N__40616\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__43428\,
            in1 => \N__40170\,
            in2 => \N__40628\,
            in3 => \N__37828\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__42966\,
            in1 => \N__40614\,
            in2 => \N__37743\,
            in3 => \N__40163\,
            lcout => \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40621\,
            in1 => \N__43319\,
            in2 => \N__40233\,
            in3 => \N__37873\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39437\,
            in2 => \N__34761\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35525\,
            in2 => \N__37443\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34737\,
            in2 => \N__35588\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35529\,
            in2 => \N__34896\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34887\,
            in2 => \N__35589\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35533\,
            in2 => \N__37515\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34881\,
            in2 => \N__35590\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35537\,
            in2 => \N__34872\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37554\,
            in2 => \N__35587\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35524\,
            in2 => \N__34860\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34848\,
            in2 => \N__35584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35512\,
            in2 => \N__37404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34917\,
            in2 => \N__35585\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35516\,
            in2 => \N__34908\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37479\,
            in2 => \N__35586\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35520\,
            in2 => \N__37347\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35414\,
            in2 => \N__37752\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37689\,
            in2 => \N__35503\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35418\,
            in2 => \N__37593\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37722\,
            in2 => \N__35504\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35422\,
            in2 => \N__37632\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34926\,
            in2 => \N__35505\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35426\,
            in2 => \N__37791\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37662\,
            in2 => \N__35506\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35401\,
            in2 => \N__37896\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_20_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37887\,
            in2 => \N__35500\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35405\,
            in2 => \N__37845\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38046\,
            in2 => \N__35501\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35409\,
            in2 => \N__37854\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38079\,
            in2 => \N__35502\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35413\,
            in2 => \N__37800\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40570\,
            in2 => \_gnd_net_\,
            in3 => \N__35301\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__35210\,
            in1 => \N__38270\,
            in2 => \_gnd_net_\,
            in3 => \N__38256\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47423\,
            ce => 'H',
            sr => \N__47062\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__35182\,
            in1 => \N__35161\,
            in2 => \_gnd_net_\,
            in3 => \N__35143\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35119\,
            in2 => \_gnd_net_\,
            in3 => \N__35098\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__35080\,
            in1 => \N__35059\,
            in2 => \N__35040\,
            in3 => \N__35035\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__35016\,
            in1 => \N__35009\,
            in2 => \N__34989\,
            in3 => \N__34985\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_14_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__36099\,
            in1 => \N__36089\,
            in2 => \N__35998\,
            in3 => \N__35846\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__38106\,
            in1 => \N__35738\,
            in2 => \N__41951\,
            in3 => \N__38214\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47549\,
            ce => 'H',
            sr => \N__46956\
        );

    \phase_controller_inst2.state_3_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__38181\,
            in1 => \N__35790\,
            in2 => \N__39583\,
            in3 => \N__38198\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47549\,
            ce => 'H',
            sr => \N__46956\
        );

    \phase_controller_inst2.T45_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35750\,
            in2 => \_gnd_net_\,
            in3 => \N__38213\,
            lcout => \T45_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47549\,
            ce => 'H',
            sr => \N__46956\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38362\,
            in2 => \_gnd_net_\,
            in3 => \N__38386\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__35739\,
            in1 => \N__41940\,
            in2 => \N__38456\,
            in3 => \N__38132\,
            lcout => \phase_controller_inst2.start_timer_tr_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_RNIG7JF_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38448\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38131\,
            lcout => \phase_controller_inst2.time_passed_RNIG7JF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36604\,
            in1 => \N__44884\,
            in2 => \_gnd_net_\,
            in3 => \N__48268\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44768\,
            in1 => \N__44201\,
            in2 => \_gnd_net_\,
            in3 => \N__48323\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47534\,
            ce => \N__47869\,
            sr => \N__46965\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44235\,
            in1 => \N__48324\,
            in2 => \_gnd_net_\,
            in3 => \N__44807\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47534\,
            ce => \N__47869\,
            sr => \N__46965\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36399\,
            in1 => \N__36459\,
            in2 => \N__44621\,
            in3 => \N__36513\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36230\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47525\,
            ce => \N__36203\,
            sr => \N__46972\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36539\,
            in1 => \N__48191\,
            in2 => \_gnd_net_\,
            in3 => \N__36514\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48190\,
            in1 => \N__36488\,
            in2 => \_gnd_net_\,
            in3 => \N__36460\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36400\,
            in1 => \N__36428\,
            in2 => \_gnd_net_\,
            in3 => \N__48192\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__36120\,
            in1 => \N__41543\,
            in2 => \N__36111\,
            in3 => \N__41522\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100001101"
        )
    port map (
            in0 => \N__41544\,
            in1 => \N__36119\,
            in2 => \N__41523\,
            in3 => \N__36107\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36663\,
            in1 => \N__48310\,
            in2 => \_gnd_net_\,
            in3 => \N__36681\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47514\,
            ce => \N__46076\,
            sr => \N__46979\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48307\,
            in1 => \N__36735\,
            in2 => \_gnd_net_\,
            in3 => \N__36756\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47514\,
            ce => \N__46076\,
            sr => \N__46979\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42283\,
            in1 => \N__48309\,
            in2 => \_gnd_net_\,
            in3 => \N__42303\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47514\,
            ce => \N__46076\,
            sr => \N__46979\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48308\,
            in1 => \N__36535\,
            in2 => \_gnd_net_\,
            in3 => \N__36515\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47514\,
            ce => \N__46076\,
            sr => \N__46979\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36484\,
            in1 => \N__36467\,
            in2 => \_gnd_net_\,
            in3 => \N__48314\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47514\,
            ce => \N__46076\,
            sr => \N__46979\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__36407\,
            in1 => \_gnd_net_\,
            in2 => \N__48339\,
            in3 => \N__36424\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47514\,
            ce => \N__46076\,
            sr => \N__46979\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__41657\,
            in1 => \N__41633\,
            in2 => \N__36267\,
            in3 => \N__36321\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__36320\,
            in1 => \N__41658\,
            in2 => \N__41637\,
            in3 => \N__36263\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36371\,
            in1 => \N__48286\,
            in2 => \_gnd_net_\,
            in3 => \N__36339\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47500\,
            ce => \N__46078\,
            sr => \N__46985\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36312\,
            in1 => \N__48322\,
            in2 => \_gnd_net_\,
            in3 => \N__36294\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47500\,
            ce => \N__46078\,
            sr => \N__46985\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44842\,
            in1 => \N__48284\,
            in2 => \_gnd_net_\,
            in3 => \N__36254\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => \elapsed_time_ns_1_RNIV8OBB_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48285\,
            in1 => \_gnd_net_\,
            in2 => \N__36618\,
            in3 => \N__44843\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47500\,
            ce => \N__46078\,
            sr => \N__46985\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36615\,
            in1 => \N__44885\,
            in2 => \_gnd_net_\,
            in3 => \N__48287\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47500\,
            ce => \N__46078\,
            sr => \N__46985\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__39113\,
            in1 => \N__36557\,
            in2 => \N__39138\,
            in3 => \N__36570\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45194\,
            in1 => \N__48247\,
            in2 => \_gnd_net_\,
            in3 => \N__45158\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => \elapsed_time_ns_1_RNIU8PBB_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48249\,
            in1 => \_gnd_net_\,
            in2 => \N__36573\,
            in3 => \N__45195\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47488\,
            ce => \N__47851\,
            sr => \N__46992\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__36569\,
            in1 => \N__39137\,
            in2 => \N__36561\,
            in3 => \N__39114\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48248\,
            in1 => \N__36540\,
            in2 => \_gnd_net_\,
            in3 => \N__36519\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47488\,
            ce => \N__47851\,
            sr => \N__46992\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36489\,
            in1 => \N__36468\,
            in2 => \_gnd_net_\,
            in3 => \N__48251\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47488\,
            ce => \N__47851\,
            sr => \N__46992\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48250\,
            in1 => \N__36429\,
            in2 => \_gnd_net_\,
            in3 => \N__36408\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47488\,
            ce => \N__47851\,
            sr => \N__46992\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41707\,
            in1 => \N__41678\,
            in2 => \_gnd_net_\,
            in3 => \N__48327\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48329\,
            in1 => \_gnd_net_\,
            in2 => \N__36765\,
            in3 => \N__41708\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47475\,
            ce => \N__47862\,
            sr => \N__47001\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36737\,
            in1 => \N__48328\,
            in2 => \_gnd_net_\,
            in3 => \N__36752\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => \elapsed_time_ns_1_RNI4EOBB_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48331\,
            in1 => \_gnd_net_\,
            in2 => \N__36741\,
            in3 => \N__36738\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47475\,
            ce => \N__47862\,
            sr => \N__47001\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__39164\,
            in1 => \N__36626\,
            in2 => \N__39189\,
            in3 => \N__36698\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__36627\,
            in1 => \N__39165\,
            in2 => \N__36702\,
            in3 => \N__39185\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36661\,
            in1 => \N__48326\,
            in2 => \_gnd_net_\,
            in3 => \N__36677\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => \elapsed_time_ns_1_RNI3DOBB_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48330\,
            in1 => \_gnd_net_\,
            in2 => \N__36666\,
            in3 => \N__36662\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47475\,
            ce => \N__47862\,
            sr => \N__47001\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46148\,
            in1 => \N__46171\,
            in2 => \_gnd_net_\,
            in3 => \N__48325\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__36983\,
            in1 => \N__46655\,
            in2 => \N__36966\,
            in3 => \N__36954\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36948\,
            in3 => \N__46558\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46559\,
            in2 => \_gnd_net_\,
            in3 => \N__36935\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39462\,
            in2 => \N__36920\,
            in3 => \N__36916\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46230\,
            in2 => \_gnd_net_\,
            in3 => \N__36852\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42507\,
            in2 => \_gnd_net_\,
            in3 => \N__36819\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42519\,
            in2 => \_gnd_net_\,
            in3 => \N__36786\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36783\,
            in2 => \_gnd_net_\,
            in3 => \N__36768\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37203\,
            in2 => \_gnd_net_\,
            in3 => \N__37167\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42543\,
            in2 => \_gnd_net_\,
            in3 => \N__37140\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42531\,
            in2 => \_gnd_net_\,
            in3 => \N__37137\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39300\,
            in2 => \_gnd_net_\,
            in3 => \N__37107\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39321\,
            in2 => \_gnd_net_\,
            in3 => \N__37080\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46335\,
            in2 => \_gnd_net_\,
            in3 => \N__37077\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42144\,
            in2 => \_gnd_net_\,
            in3 => \N__37041\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42153\,
            in2 => \_gnd_net_\,
            in3 => \N__36999\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36996\,
            in2 => \_gnd_net_\,
            in3 => \N__36987\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39639\,
            in2 => \_gnd_net_\,
            in3 => \N__37257\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39621\,
            in2 => \_gnd_net_\,
            in3 => \N__37254\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39306\,
            in2 => \_gnd_net_\,
            in3 => \N__37251\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_15_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39612\,
            in2 => \_gnd_net_\,
            in3 => \N__37248\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39312\,
            in2 => \_gnd_net_\,
            in3 => \N__37245\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39327\,
            in2 => \_gnd_net_\,
            in3 => \N__37242\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39645\,
            in2 => \_gnd_net_\,
            in3 => \N__37212\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46188\,
            in2 => \_gnd_net_\,
            in3 => \N__37209\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46287\,
            in2 => \_gnd_net_\,
            in3 => \N__37206\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39630\,
            in2 => \_gnd_net_\,
            in3 => \N__37308\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37506\,
            in2 => \_gnd_net_\,
            in3 => \N__37305\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_15_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39516\,
            in2 => \_gnd_net_\,
            in3 => \N__37302\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39507\,
            in2 => \_gnd_net_\,
            in3 => \N__37299\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42135\,
            in2 => \_gnd_net_\,
            in3 => \N__37296\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41316\,
            in2 => \_gnd_net_\,
            in3 => \N__37293\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37290\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110110001"
        )
    port map (
            in0 => \N__40594\,
            in1 => \N__42932\,
            in2 => \N__37656\,
            in3 => \N__40175\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__40174\,
            in1 => \N__40595\,
            in2 => \N__46323\,
            in3 => \N__37682\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42400\,
            in1 => \N__38012\,
            in2 => \_gnd_net_\,
            in3 => \N__37537\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43416\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42581\,
            in1 => \N__38014\,
            in2 => \_gnd_net_\,
            in3 => \N__37499\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__38011\,
            in1 => \N__37471\,
            in2 => \_gnd_net_\,
            in3 => \N__39490\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46372\,
            in1 => \N__38013\,
            in2 => \_gnd_net_\,
            in3 => \N__37423\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40581\,
            in1 => \N__43391\,
            in2 => \N__40266\,
            in3 => \N__40291\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__43132\,
            in1 => \N__37372\,
            in2 => \_gnd_net_\,
            in3 => \N__38015\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__40228\,
            in1 => \N__40582\,
            in2 => \N__39452\,
            in3 => \N__39406\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40625\,
            in1 => \N__43473\,
            in2 => \N__40267\,
            in3 => \N__37917\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__39365\,
            in1 => \N__46217\,
            in2 => \_gnd_net_\,
            in3 => \N__38039\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38034\,
            in1 => \N__43087\,
            in2 => \_gnd_net_\,
            in3 => \N__37775\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__37742\,
            in1 => \N__38037\,
            in2 => \_gnd_net_\,
            in3 => \N__42959\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38035\,
            in1 => \N__43046\,
            in2 => \_gnd_net_\,
            in3 => \N__37712\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__46318\,
            in1 => \N__37683\,
            in2 => \_gnd_net_\,
            in3 => \N__38040\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38038\,
            in1 => \N__42931\,
            in2 => \_gnd_net_\,
            in3 => \N__37655\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__42997\,
            in1 => \N__37616\,
            in2 => \_gnd_net_\,
            in3 => \N__38036\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38017\,
            in1 => \N__42796\,
            in2 => \_gnd_net_\,
            in3 => \N__37574\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40611\,
            in1 => \N__46218\,
            in2 => \N__40268\,
            in3 => \N__39369\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43273\,
            in1 => \N__40610\,
            in2 => \_gnd_net_\,
            in3 => \N__38314\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40608\,
            in1 => \N__43346\,
            in2 => \_gnd_net_\,
            in3 => \N__38063\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__38018\,
            in1 => \N__43471\,
            in2 => \_gnd_net_\,
            in3 => \N__37916\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40606\,
            in1 => \N__43426\,
            in2 => \_gnd_net_\,
            in3 => \N__37829\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43312\,
            in1 => \N__40609\,
            in2 => \_gnd_net_\,
            in3 => \N__37874\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40607\,
            in1 => \N__43390\,
            in2 => \_gnd_net_\,
            in3 => \N__40293\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__40246\,
            in1 => \N__40565\,
            in2 => \N__37836\,
            in3 => \N__43427\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40564\,
            in2 => \_gnd_net_\,
            in3 => \N__39411\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__40566\,
            in1 => \N__40245\,
            in2 => \N__43280\,
            in3 => \N__38316\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_tr_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38248\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38226\,
            ce => 'H',
            sr => \N__47063\
        );

    \delay_measurement_inst.start_timer_tr_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38247\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38225\,
            ce => 'H',
            sr => \N__47064\
        );

    \phase_controller_inst2.state_RNI9M3O_0_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38104\,
            in2 => \_gnd_net_\,
            in3 => \N__38212\,
            lcout => \phase_controller_inst2.state_RNI9M3OZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46957\
        );

    \phase_controller_inst2.stoper_tr.running_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000011111100"
        )
    port map (
            in0 => \N__38882\,
            in1 => \N__41283\,
            in2 => \N__38406\,
            in3 => \N__38366\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46957\
        );

    \phase_controller_inst2.start_timer_tr_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__38199\,
            in1 => \N__38187\,
            in2 => \N__38391\,
            in3 => \N__46467\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46957\
        );

    \phase_controller_inst2.state_2_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__38173\,
            in1 => \N__38133\,
            in2 => \N__38457\,
            in3 => \N__39575\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46957\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010100100000"
        )
    port map (
            in0 => \N__41282\,
            in1 => \N__38883\,
            in2 => \N__38367\,
            in3 => \N__38105\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46957\
        );

    \phase_controller_inst2.T12_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__38455\,
            in1 => \N__38417\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \T12_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47550\,
            ce => 'H',
            sr => \N__46957\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__38402\,
            in1 => \N__38361\,
            in2 => \_gnd_net_\,
            in3 => \N__38385\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41279\,
            in2 => \_gnd_net_\,
            in3 => \N__41258\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101011101"
        )
    port map (
            in0 => \N__38360\,
            in1 => \N__41871\,
            in2 => \N__41853\,
            in3 => \N__38898\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38340\,
            in3 => \N__41280\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__41495\,
            in1 => \N__41471\,
            in2 => \N__38328\,
            in3 => \N__38337\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__38336\,
            in1 => \N__41496\,
            in2 => \N__41475\,
            in3 => \N__38324\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45279\,
            in1 => \N__45316\,
            in2 => \_gnd_net_\,
            in3 => \N__48228\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47535\,
            ce => \N__46077\,
            sr => \N__46966\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48225\,
            in1 => \N__44259\,
            in2 => \_gnd_net_\,
            in3 => \N__44298\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47535\,
            ce => \N__46077\,
            sr => \N__46966\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44617\,
            in1 => \N__44643\,
            in2 => \_gnd_net_\,
            in3 => \N__48229\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47535\,
            ce => \N__46077\,
            sr => \N__46966\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48226\,
            in1 => \N__44767\,
            in2 => \_gnd_net_\,
            in3 => \N__44205\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47535\,
            ce => \N__46077\,
            sr => \N__46966\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44805\,
            in1 => \N__44234\,
            in2 => \_gnd_net_\,
            in3 => \N__48230\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47535\,
            ce => \N__46077\,
            sr => \N__46966\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48227\,
            in1 => \N__45345\,
            in2 => \_gnd_net_\,
            in3 => \N__45370\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47535\,
            ce => \N__46077\,
            sr => \N__46966\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40715\,
            in1 => \N__38538\,
            in2 => \N__38532\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38523\,
            in2 => \N__38514\,
            in3 => \N__40682\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38505\,
            in2 => \N__38496\,
            in3 => \N__40658\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40643\,
            in1 => \N__38487\,
            in2 => \N__38481\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38463\,
            in2 => \N__38472\,
            in3 => \N__41444\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38637\,
            in2 => \N__38631\,
            in3 => \N__41430\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38622\,
            in2 => \N__38616\,
            in3 => \N__41408\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46095\,
            in2 => \N__38604\,
            in3 => \N__41393\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41379\,
            in1 => \N__38595\,
            in2 => \N__45027\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44952\,
            in2 => \N__38589\,
            in3 => \N__41360\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41345\,
            in1 => \N__38580\,
            in2 => \N__38574\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38565\,
            in2 => \N__38559\,
            in3 => \N__41330\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46107\,
            in2 => \N__38550\,
            in3 => \N__41588\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41573\,
            in1 => \N__41667\,
            in2 => \N__38715\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__41558\,
            in1 => \N__38697\,
            in2 => \N__38706\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38691\,
            in2 => \N__38685\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38676\,
            in2 => \N__38667\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45255\,
            in2 => \N__45210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38652\,
            in2 => \N__38646\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44940\,
            in2 => \N__44898\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45504\,
            in2 => \N__45453\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45441\,
            in2 => \N__45393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41867\,
            in2 => \N__41733\,
            in3 => \N__38889\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38886\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38868\,
            in2 => \N__38862\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47837\,
            in1 => \N__38822\,
            in2 => \_gnd_net_\,
            in3 => \N__38808\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__47841\,
            in1 => \N__38789\,
            in2 => \N__38805\,
            in3 => \N__38775\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47838\,
            in1 => \N__38771\,
            in2 => \_gnd_net_\,
            in3 => \N__38757\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47842\,
            in1 => \N__38753\,
            in2 => \_gnd_net_\,
            in3 => \N__38739\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47839\,
            in1 => \N__38732\,
            in2 => \_gnd_net_\,
            in3 => \N__38718\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47843\,
            in1 => \N__39041\,
            in2 => \_gnd_net_\,
            in3 => \N__39027\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47840\,
            in1 => \N__39023\,
            in2 => \_gnd_net_\,
            in3 => \N__39009\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__47489\,
            ce => 'H',
            sr => \N__46993\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47850\,
            in1 => \N__39005\,
            in2 => \_gnd_net_\,
            in3 => \N__38991\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47777\,
            in1 => \N__38987\,
            in2 => \_gnd_net_\,
            in3 => \N__38973\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47847\,
            in1 => \N__38969\,
            in2 => \_gnd_net_\,
            in3 => \N__38955\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47778\,
            in1 => \N__38951\,
            in2 => \_gnd_net_\,
            in3 => \N__38937\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47848\,
            in1 => \N__38933\,
            in2 => \_gnd_net_\,
            in3 => \N__38919\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47779\,
            in1 => \N__38915\,
            in2 => \_gnd_net_\,
            in3 => \N__38901\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47849\,
            in1 => \N__39206\,
            in2 => \_gnd_net_\,
            in3 => \N__39192\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47780\,
            in1 => \N__39184\,
            in2 => \_gnd_net_\,
            in3 => \N__39168\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__47476\,
            ce => 'H',
            sr => \N__47002\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47833\,
            in1 => \N__39163\,
            in2 => \_gnd_net_\,
            in3 => \N__39147\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47819\,
            in1 => \N__42231\,
            in2 => \_gnd_net_\,
            in3 => \N__39144\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47834\,
            in1 => \N__42192\,
            in2 => \_gnd_net_\,
            in3 => \N__39141\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47820\,
            in1 => \N__39133\,
            in2 => \_gnd_net_\,
            in3 => \N__39117\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47835\,
            in1 => \N__39112\,
            in2 => \_gnd_net_\,
            in3 => \N__39096\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47821\,
            in1 => \N__39083\,
            in2 => \_gnd_net_\,
            in3 => \N__39069\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47836\,
            in1 => \N__39059\,
            in2 => \_gnd_net_\,
            in3 => \N__39045\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47822\,
            in1 => \N__45854\,
            in2 => \_gnd_net_\,
            in3 => \N__39291\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__47464\,
            ce => 'H',
            sr => \N__47008\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47829\,
            in1 => \N__45839\,
            in2 => \_gnd_net_\,
            in3 => \N__39288\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_16_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47826\,
            in1 => \N__45926\,
            in2 => \_gnd_net_\,
            in3 => \N__39285\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47830\,
            in1 => \N__45953\,
            in2 => \_gnd_net_\,
            in3 => \N__39282\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47827\,
            in1 => \N__46037\,
            in2 => \_gnd_net_\,
            in3 => \N__39279\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47831\,
            in1 => \N__46013\,
            in2 => \_gnd_net_\,
            in3 => \N__39276\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47828\,
            in1 => \N__39257\,
            in2 => \_gnd_net_\,
            in3 => \N__39243\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__47832\,
            in1 => \N__39224\,
            in2 => \_gnd_net_\,
            in3 => \N__39240\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47456\,
            ce => 'H',
            sr => \N__47014\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43710\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47446\,
            ce => \N__43231\,
            sr => \N__47021\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39480\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \N__39453\,
            in1 => \N__40629\,
            in2 => \N__40271\,
            in3 => \N__39407\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__40596\,
            in1 => \N__46210\,
            in2 => \N__40269\,
            in3 => \N__39364\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42913\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42694\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42947\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43029\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42732\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__40597\,
            in1 => \N__40292\,
            in2 => \N__40270\,
            in3 => \N__43392\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42874\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43114\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43452\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43069\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42980\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.T01_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39527\,
            in2 => \_gnd_net_\,
            in3 => \N__39599\,
            lcout => \T01_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47435\,
            ce => 'H',
            sr => \N__47033\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43372\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43334\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43254\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41307\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44251\,
            in1 => \N__44297\,
            in2 => \_gnd_net_\,
            in3 => \N__48189\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47554\,
            ce => \N__47824\,
            sr => \N__46955\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__41281\,
            in1 => \N__41259\,
            in2 => \N__40716\,
            in3 => \N__42122\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47551\,
            ce => 'H',
            sr => \N__46958\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40738\,
            in1 => \N__41247\,
            in2 => \_gnd_net_\,
            in3 => \N__41186\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40711\,
            in2 => \N__40692\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42092\,
            in1 => \N__40683\,
            in2 => \_gnd_net_\,
            in3 => \N__40671\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__42096\,
            in1 => \N__40668\,
            in2 => \N__40662\,
            in3 => \N__40647\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42093\,
            in1 => \N__40644\,
            in2 => \_gnd_net_\,
            in3 => \N__40632\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42097\,
            in1 => \N__41445\,
            in2 => \_gnd_net_\,
            in3 => \N__41433\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42094\,
            in1 => \N__41426\,
            in2 => \_gnd_net_\,
            in3 => \N__41412\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42098\,
            in1 => \N__41409\,
            in2 => \_gnd_net_\,
            in3 => \N__41397\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42095\,
            in1 => \N__41394\,
            in2 => \_gnd_net_\,
            in3 => \N__41382\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__47545\,
            ce => 'H',
            sr => \N__46961\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42106\,
            in1 => \N__41378\,
            in2 => \_gnd_net_\,
            in3 => \N__41364\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42099\,
            in1 => \N__41361\,
            in2 => \_gnd_net_\,
            in3 => \N__41349\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42103\,
            in1 => \N__41346\,
            in2 => \_gnd_net_\,
            in3 => \N__41334\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42100\,
            in1 => \N__41331\,
            in2 => \_gnd_net_\,
            in3 => \N__41319\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42104\,
            in1 => \N__41589\,
            in2 => \_gnd_net_\,
            in3 => \N__41577\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42101\,
            in1 => \N__41574\,
            in2 => \_gnd_net_\,
            in3 => \N__41562\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42105\,
            in1 => \N__41559\,
            in2 => \_gnd_net_\,
            in3 => \N__41547\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42102\,
            in1 => \N__41542\,
            in2 => \_gnd_net_\,
            in3 => \N__41526\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__47536\,
            ce => 'H',
            sr => \N__46967\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42107\,
            in1 => \N__41513\,
            in2 => \_gnd_net_\,
            in3 => \N__41499\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42111\,
            in1 => \N__41494\,
            in2 => \_gnd_net_\,
            in3 => \N__41478\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42108\,
            in1 => \N__41470\,
            in2 => \_gnd_net_\,
            in3 => \N__41454\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42112\,
            in1 => \N__45227\,
            in2 => \_gnd_net_\,
            in3 => \N__41451\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42109\,
            in1 => \N__45243\,
            in2 => \_gnd_net_\,
            in3 => \N__41448\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42113\,
            in1 => \N__41656\,
            in2 => \_gnd_net_\,
            in3 => \N__41640\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42110\,
            in1 => \N__41632\,
            in2 => \_gnd_net_\,
            in3 => \N__41613\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42114\,
            in1 => \N__44915\,
            in2 => \_gnd_net_\,
            in3 => \N__41610\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__47526\,
            ce => 'H',
            sr => \N__46973\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42115\,
            in1 => \N__44931\,
            in2 => \_gnd_net_\,
            in3 => \N__41607\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42119\,
            in1 => \N__45479\,
            in2 => \_gnd_net_\,
            in3 => \N__41604\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42116\,
            in1 => \N__45495\,
            in2 => \_gnd_net_\,
            in3 => \N__41601\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42120\,
            in1 => \N__45428\,
            in2 => \_gnd_net_\,
            in3 => \N__41598\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42117\,
            in1 => \N__45410\,
            in2 => \_gnd_net_\,
            in3 => \N__41595\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42121\,
            in1 => \N__41755\,
            in2 => \_gnd_net_\,
            in3 => \N__41592\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__42118\,
            in1 => \N__41775\,
            in2 => \_gnd_net_\,
            in3 => \N__41958\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.T23_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41882\,
            in2 => \_gnd_net_\,
            in3 => \N__41944\,
            lcout => \T23_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47515\,
            ce => 'H',
            sr => \N__46980\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100001010"
        )
    port map (
            in0 => \N__41772\,
            in1 => \N__41748\,
            in2 => \N__41724\,
            in3 => \N__41786\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__41785\,
            in1 => \N__41773\,
            in2 => \N__41756\,
            in3 => \N__41719\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_df30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48340\,
            in1 => \N__41838\,
            in2 => \_gnd_net_\,
            in3 => \N__41805\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47501\,
            ce => \N__46080\,
            sr => \N__46986\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__41787\,
            in1 => \N__41774\,
            in2 => \N__41757\,
            in3 => \N__41723\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48341\,
            in1 => \N__44716\,
            in2 => \_gnd_net_\,
            in3 => \N__44325\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47501\,
            ce => \N__46080\,
            sr => \N__46986\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41709\,
            in1 => \N__41682\,
            in2 => \_gnd_net_\,
            in3 => \N__48342\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47501\,
            ce => \N__46080\,
            sr => \N__46986\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__42242\,
            in1 => \N__42190\,
            in2 => \N__42212\,
            in3 => \N__42229\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42284\,
            in1 => \N__48294\,
            in2 => \_gnd_net_\,
            in3 => \N__42296\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => \elapsed_time_ns_1_RNI2COBB_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__48295\,
            in1 => \N__42285\,
            in2 => \N__42255\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47490\,
            ce => \N__47815\,
            sr => \N__46994\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45318\,
            in1 => \N__45271\,
            in2 => \_gnd_net_\,
            in3 => \N__48296\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47490\,
            ce => \N__47815\,
            sr => \N__46994\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110010"
        )
    port map (
            in0 => \N__42243\,
            in1 => \N__42230\,
            in2 => \N__42213\,
            in3 => \N__42191\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__45905\,
            in1 => \N__45949\,
            in2 => \N__45978\,
            in3 => \N__45925\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42604\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42651\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__43303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42820\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42777\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42427\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42472\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43166\,
            in2 => \N__43679\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43706\,
            in2 => \N__43650\,
            in3 => \N__42456\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43680\,
            in2 => \N__43619\,
            in3 => \N__42411\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43649\,
            in2 => \N__43589\,
            in3 => \N__42363\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43559\,
            in2 => \N__43620\,
            in3 => \N__42321\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43532\,
            in2 => \N__43590\,
            in3 => \N__42804\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43560\,
            in2 => \N__43505\,
            in3 => \N__42759\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43955\,
            in2 => \N__43536\,
            in3 => \N__42717\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__47457\,
            ce => \N__43233\,
            sr => \N__47015\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43928\,
            in2 => \N__43506\,
            in3 => \N__42678\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43907\,
            in2 => \N__43962\,
            in3 => \N__42675\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43929\,
            in2 => \N__43884\,
            in3 => \N__42624\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43908\,
            in2 => \N__43856\,
            in3 => \N__42585\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43883\,
            in2 => \N__43826\,
            in3 => \N__42546\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43796\,
            in2 => \N__43857\,
            in3 => \N__43098\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43769\,
            in2 => \N__43827\,
            in3 => \N__43053\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43797\,
            in2 => \N__43743\,
            in3 => \N__43011\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__47447\,
            ce => \N__43232\,
            sr => \N__47022\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44174\,
            in2 => \N__43773\,
            in3 => \N__42969\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43742\,
            in2 => \N__44147\,
            in3 => \N__42936\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44120\,
            in2 => \N__44178\,
            in3 => \N__42897\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44096\,
            in2 => \N__44148\,
            in3 => \N__42861\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44121\,
            in2 => \N__44072\,
            in3 => \N__42858\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44045\,
            in2 => \N__44100\,
            in3 => \N__42855\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44021\,
            in2 => \N__44073\,
            in3 => \N__43431\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44046\,
            in2 => \N__43994\,
            in3 => \N__43395\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__47441\,
            ce => \N__43230\,
            sr => \N__47028\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44570\,
            in2 => \N__44025\,
            in3 => \N__43356\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__47436\,
            ce => \N__43228\,
            sr => \N__47034\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43995\,
            in2 => \N__44543\,
            in3 => \N__43323\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__47436\,
            ce => \N__43228\,
            sr => \N__47034\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44517\,
            in2 => \N__44574\,
            in3 => \N__43284\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__47436\,
            ce => \N__43228\,
            sr => \N__47034\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44379\,
            in2 => \N__44544\,
            in3 => \N__43236\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__47436\,
            ce => \N__43228\,
            sr => \N__47034\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43203\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44489\,
            in1 => \N__43162\,
            in2 => \_gnd_net_\,
            in3 => \N__43143\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_1_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44485\,
            in1 => \N__43702\,
            in2 => \_gnd_net_\,
            in3 => \N__43683\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_2_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44490\,
            in1 => \N__43672\,
            in2 => \_gnd_net_\,
            in3 => \N__43653\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_3_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44486\,
            in1 => \N__43639\,
            in2 => \_gnd_net_\,
            in3 => \N__43623\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_4_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44491\,
            in1 => \N__43607\,
            in2 => \_gnd_net_\,
            in3 => \N__43593\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_5_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44487\,
            in1 => \N__43577\,
            in2 => \_gnd_net_\,
            in3 => \N__43563\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_6_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44492\,
            in1 => \N__43553\,
            in2 => \_gnd_net_\,
            in3 => \N__43539\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_7_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44488\,
            in1 => \N__43525\,
            in2 => \_gnd_net_\,
            in3 => \N__43509\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__47432\,
            ce => \N__44356\,
            sr => \N__47040\
        );

    \current_shift_inst.timer_s1.counter_8_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44496\,
            in1 => \N__43492\,
            in2 => \_gnd_net_\,
            in3 => \N__43476\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_9_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44477\,
            in1 => \N__43954\,
            in2 => \_gnd_net_\,
            in3 => \N__43932\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_10_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44493\,
            in1 => \N__43927\,
            in2 => \_gnd_net_\,
            in3 => \N__43911\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_11_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44474\,
            in1 => \N__43901\,
            in2 => \_gnd_net_\,
            in3 => \N__43887\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_12_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44494\,
            in1 => \N__43879\,
            in2 => \_gnd_net_\,
            in3 => \N__43860\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_13_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44475\,
            in1 => \N__43844\,
            in2 => \_gnd_net_\,
            in3 => \N__43830\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_14_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44495\,
            in1 => \N__43814\,
            in2 => \_gnd_net_\,
            in3 => \N__43800\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_15_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44476\,
            in1 => \N__43790\,
            in2 => \_gnd_net_\,
            in3 => \N__43776\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__47428\,
            ce => \N__44363\,
            sr => \N__47045\
        );

    \current_shift_inst.timer_s1.counter_16_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44470\,
            in1 => \N__43762\,
            in2 => \_gnd_net_\,
            in3 => \N__43746\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_17_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44481\,
            in1 => \N__43732\,
            in2 => \_gnd_net_\,
            in3 => \N__43713\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_18_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44471\,
            in1 => \N__44167\,
            in2 => \_gnd_net_\,
            in3 => \N__44151\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_19_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44482\,
            in1 => \N__44140\,
            in2 => \_gnd_net_\,
            in3 => \N__44124\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_20_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44472\,
            in1 => \N__44119\,
            in2 => \_gnd_net_\,
            in3 => \N__44103\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_21_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44483\,
            in1 => \N__44095\,
            in2 => \_gnd_net_\,
            in3 => \N__44076\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_22_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44473\,
            in1 => \N__44065\,
            in2 => \_gnd_net_\,
            in3 => \N__44049\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_23_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44484\,
            in1 => \N__44044\,
            in2 => \_gnd_net_\,
            in3 => \N__44028\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__47427\,
            ce => \N__44355\,
            sr => \N__47051\
        );

    \current_shift_inst.timer_s1.counter_24_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44497\,
            in1 => \N__44014\,
            in2 => \_gnd_net_\,
            in3 => \N__43998\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__47426\,
            ce => \N__44364\,
            sr => \N__47055\
        );

    \current_shift_inst.timer_s1.counter_25_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44478\,
            in1 => \N__43987\,
            in2 => \_gnd_net_\,
            in3 => \N__43965\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__47426\,
            ce => \N__44364\,
            sr => \N__47055\
        );

    \current_shift_inst.timer_s1.counter_26_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44498\,
            in1 => \N__44563\,
            in2 => \_gnd_net_\,
            in3 => \N__44547\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__47426\,
            ce => \N__44364\,
            sr => \N__47055\
        );

    \current_shift_inst.timer_s1.counter_27_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44479\,
            in1 => \N__44536\,
            in2 => \_gnd_net_\,
            in3 => \N__44520\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__47426\,
            ce => \N__44364\,
            sr => \N__47055\
        );

    \current_shift_inst.timer_s1.counter_28_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44499\,
            in1 => \N__44516\,
            in2 => \_gnd_net_\,
            in3 => \N__44502\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__47426\,
            ce => \N__44364\,
            sr => \N__47055\
        );

    \current_shift_inst.timer_s1.counter_29_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44480\,
            in1 => \N__44378\,
            in2 => \_gnd_net_\,
            in3 => \N__44382\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47426\,
            ce => \N__44364\,
            sr => \N__47055\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44320\,
            in1 => \N__44721\,
            in2 => \_gnd_net_\,
            in3 => \N__48188\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48187\,
            in1 => \N__44255\,
            in2 => \_gnd_net_\,
            in3 => \N__44296\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48042\,
            in1 => \N__44808\,
            in2 => \_gnd_net_\,
            in3 => \N__44233\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_18_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44200\,
            in1 => \N__44769\,
            in2 => \_gnd_net_\,
            in3 => \N__48043\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_18_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48041\,
            in1 => \N__45010\,
            in2 => \_gnd_net_\,
            in3 => \N__44990\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48448\,
            in2 => \_gnd_net_\,
            in3 => \N__45369\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__44886\,
            in1 => \N__44976\,
            in2 => \N__44847\,
            in3 => \N__45051\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__44806\,
            in1 => \N__44754\,
            in2 => \N__44730\,
            in3 => \N__44727\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__44717\,
            in1 => \N__44676\,
            in2 => \N__44664\,
            in3 => \N__44649\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__45052\,
            in1 => \_gnd_net_\,
            in2 => \N__44661\,
            in3 => \N__45079\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__45586\,
            in1 => \N__45648\,
            in2 => \_gnd_net_\,
            in3 => \N__44658\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44642\,
            in1 => \N__44616\,
            in2 => \_gnd_net_\,
            in3 => \N__48044\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45543\,
            in1 => \N__48073\,
            in2 => \_gnd_net_\,
            in3 => \N__45561\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47546\,
            ce => \N__47873\,
            sr => \N__46962\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44638\,
            in1 => \N__44622\,
            in2 => \_gnd_net_\,
            in3 => \N__48074\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47546\,
            ce => \N__47873\,
            sr => \N__46962\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__45242\,
            in1 => \N__45223\,
            in2 => \N__45096\,
            in3 => \N__45147\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__45146\,
            in1 => \N__45241\,
            in2 => \N__45228\,
            in3 => \N__45092\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__48184\,
            in1 => \N__45193\,
            in2 => \_gnd_net_\,
            in3 => \N__45165\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47537\,
            ce => \N__46079\,
            sr => \N__46968\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45138\,
            in1 => \N__48186\,
            in2 => \_gnd_net_\,
            in3 => \N__45117\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47537\,
            ce => \N__46079\,
            sr => \N__46968\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48185\,
            in1 => \N__45080\,
            in2 => \_gnd_net_\,
            in3 => \N__45060\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47537\,
            ce => \N__46079\,
            sr => \N__46968\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45011\,
            in1 => \N__44991\,
            in2 => \_gnd_net_\,
            in3 => \N__48120\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47537\,
            ce => \N__46079\,
            sr => \N__46968\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__44930\,
            in1 => \N__45677\,
            in2 => \N__44916\,
            in3 => \N__45708\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__45707\,
            in1 => \N__44929\,
            in2 => \N__45681\,
            in3 => \N__44914\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45541\,
            in1 => \N__48118\,
            in2 => \_gnd_net_\,
            in3 => \N__45557\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => \elapsed_time_ns_1_RNI4FPBB_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48119\,
            in1 => \_gnd_net_\,
            in2 => \N__45546\,
            in3 => \N__45542\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47527\,
            ce => \N__46081\,
            sr => \N__46974\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__45461\,
            in1 => \N__45478\,
            in2 => \N__45696\,
            in3 => \N__45493\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__45494\,
            in1 => \N__45692\,
            in2 => \N__45480\,
            in3 => \N__45462\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__45717\,
            in1 => \N__45726\,
            in2 => \N__45429\,
            in3 => \N__45409\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__45725\,
            in1 => \N__45427\,
            in2 => \N__45411\,
            in3 => \N__45716\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48257\,
            in1 => \N__45344\,
            in2 => \_gnd_net_\,
            in3 => \N__45377\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45275\,
            in1 => \N__45317\,
            in2 => \_gnd_net_\,
            in3 => \N__48256\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45597\,
            in1 => \N__48301\,
            in2 => \_gnd_net_\,
            in3 => \N__45612\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47502\,
            ce => \N__46083\,
            sr => \N__46987\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48298\,
            in1 => \N__48405\,
            in2 => \_gnd_net_\,
            in3 => \N__48377\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47502\,
            ce => \N__46083\,
            sr => \N__46987\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46509\,
            in1 => \N__48299\,
            in2 => \_gnd_net_\,
            in3 => \N__45741\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47502\,
            ce => \N__46083\,
            sr => \N__46987\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__48297\,
            in1 => \N__45666\,
            in2 => \_gnd_net_\,
            in3 => \N__45651\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47502\,
            ce => \N__46083\,
            sr => \N__46987\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45786\,
            in1 => \N__48300\,
            in2 => \_gnd_net_\,
            in3 => \N__45804\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47502\,
            ce => \N__46083\,
            sr => \N__46987\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45649\,
            in1 => \N__48258\,
            in2 => \_gnd_net_\,
            in3 => \N__45665\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48260\,
            in1 => \_gnd_net_\,
            in2 => \N__45654\,
            in3 => \N__45650\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47491\,
            ce => \N__47811\,
            sr => \N__46995\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45595\,
            in1 => \N__48259\,
            in2 => \_gnd_net_\,
            in3 => \N__45611\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => \elapsed_time_ns_1_RNI6HPBB_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48261\,
            in1 => \_gnd_net_\,
            in2 => \N__45600\,
            in3 => \N__45596\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47491\,
            ce => \N__47811\,
            sr => \N__46995\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__45998\,
            in1 => \N__46044\,
            in2 => \N__46023\,
            in3 => \N__47891\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__46043\,
            in1 => \N__46022\,
            in2 => \N__47895\,
            in3 => \N__45999\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000010"
        )
    port map (
            in0 => \N__45977\,
            in1 => \N__45957\,
            in2 => \N__45933\,
            in3 => \N__45906\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__45750\,
            in1 => \N__46476\,
            in2 => \N__45864\,
            in3 => \N__45835\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__46475\,
            in1 => \N__45863\,
            in2 => \N__45840\,
            in3 => \N__45749\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45781\,
            in1 => \N__48253\,
            in2 => \_gnd_net_\,
            in3 => \N__45800\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48255\,
            in1 => \_gnd_net_\,
            in2 => \N__45789\,
            in3 => \N__45782\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47477\,
            ce => \N__47823\,
            sr => \N__47003\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46501\,
            in1 => \N__48252\,
            in2 => \_gnd_net_\,
            in3 => \N__45737\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => \elapsed_time_ns_1_RNI2DPBB_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__48254\,
            in1 => \_gnd_net_\,
            in2 => \N__46512\,
            in3 => \N__46502\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47477\,
            ce => \N__47823\,
            sr => \N__47003\
        );

    \phase_controller_inst1.start_timer_tr_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__46455\,
            in1 => \N__46413\,
            in2 => \N__46592\,
            in3 => \N__46398\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47465\,
            ce => 'H',
            sr => \N__47009\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__46587\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47465\,
            ce => 'H',
            sr => \N__47009\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46353\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46300\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46248\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46204\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46176\,
            in1 => \N__46152\,
            in2 => \_gnd_net_\,
            in3 => \N__48305\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47555\,
            ce => \N__46082\,
            sr => \N__46963\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48421\,
            in1 => \N__48465\,
            in2 => \_gnd_net_\,
            in3 => \N__48306\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47555\,
            ce => \N__46082\,
            sr => \N__46963\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48425\,
            in1 => \N__48464\,
            in2 => \_gnd_net_\,
            in3 => \N__48293\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48400\,
            in1 => \N__48376\,
            in2 => \_gnd_net_\,
            in3 => \N__48262\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48401\,
            in1 => \N__48378\,
            in2 => \_gnd_net_\,
            in3 => \N__48338\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47528\,
            ce => \N__47735\,
            sr => \N__46988\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46650\,
            in2 => \_gnd_net_\,
            in3 => \N__46593\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111110000"
        )
    port map (
            in0 => \N__46651\,
            in1 => \N__47583\,
            in2 => \N__46608\,
            in3 => \N__46536\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47503\,
            ce => 'H',
            sr => \N__47004\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__46637\,
            in1 => \N__46604\,
            in2 => \_gnd_net_\,
            in3 => \N__46588\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
