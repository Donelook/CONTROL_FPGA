-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 8 2025 23:57:57

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    start_stop : in std_logic;
    s2_phy : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__22544\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22238\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22051\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17291\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \bfn_1_18_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \bfn_1_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_1_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \N_27_i_i\ : std_logic;
signal un7_start_stop : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_2_17_0_\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \bfn_2_22_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\ : std_logic;
signal \bfn_2_23_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \delay_measurement_inst.N_212_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_3_21_0_\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \delay_measurement_inst.N_168\ : std_logic;
signal \delay_measurement_inst.N_81_i\ : std_logic;
signal \delay_measurement_inst.N_81_i_cascade_\ : std_logic;
signal \delay_measurement_inst.N_200\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\ : std_logic;
signal \delay_measurement_inst.un1_tr_state_1_i_0_a2_0_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_203\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_3\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_11\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_4_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \bfn_4_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_138_i_g\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_slave.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_15_cascade_\ : std_logic;
signal il_max_comp2_c : std_logic;
signal \il_max_comp2_D1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6Z0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_92_cascade_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\ : std_logic;
signal \delay_measurement_inst.N_165\ : std_logic;
signal \delay_measurement_inst.N_212\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_18\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_19\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\ : std_logic;
signal \delay_measurement_inst.N_197_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.N_81_i_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_5_17_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_5_18_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_139_i_g\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m3_eZ0Z_1\ : std_logic;
signal phase_controller_inst1_stoper_hc_un1_startlto19_2 : std_logic;
signal \phase_controller_inst1_stoper_hc_un1_startlto19_2_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_a0Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_aZ0Z2_cascade_\ : std_logic;
signal \d_N_5_mux\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_2_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_N_6_mux\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_m2_eZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal measured_delay_tr_11 : std_logic;
signal measured_delay_tr_9 : std_logic;
signal \phase_controller_inst1.stoper_tr.N_98\ : std_logic;
signal measured_delay_tr_12 : std_logic;
signal measured_delay_tr_13 : std_logic;
signal measured_delay_tr_14 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\ : std_logic;
signal measured_delay_tr_10 : std_logic;
signal measured_delay_tr_4 : std_logic;
signal measured_delay_tr_7 : std_logic;
signal measured_delay_tr_8 : std_logic;
signal measured_delay_tr_5 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\ : std_logic;
signal measured_delay_tr_1 : std_logic;
signal measured_delay_tr_2 : std_logic;
signal measured_delay_tr_3 : std_logic;
signal \phase_controller_inst1.stoper_tr.N_109\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_110\ : std_logic;
signal \phase_controller_inst1.stoper_tr.N_92\ : std_logic;
signal measured_delay_tr_6 : std_logic;
signal \phase_controller_inst1.stoper_tr.N_95\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_17\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal measured_delay_tr_19 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal measured_delay_tr_17 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal measured_delay_tr_18 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal measured_delay_tr_16 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlt31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_16\ : std_logic;
signal \bfn_7_21_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal measured_delay_hc_4 : std_logic;
signal measured_delay_hc_1 : std_logic;
signal measured_delay_hc_22 : std_logic;
signal measured_delay_hc_21 : std_logic;
signal measured_delay_hc_0 : std_logic;
signal measured_delay_hc_5 : std_logic;
signal measured_delay_hc_20 : std_logic;
signal measured_delay_hc_3 : std_logic;
signal measured_delay_hc_17 : std_logic;
signal measured_delay_hc_6 : std_logic;
signal measured_delay_hc_13 : std_logic;
signal measured_delay_hc_19 : std_logic;
signal measured_delay_hc_15 : std_logic;
signal measured_delay_hc_18 : std_logic;
signal measured_delay_hc_16 : std_logic;
signal measured_delay_hc_14 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\ : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11_cascade_\ : std_logic;
signal \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_slave.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_start\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_startlto31_d\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal measured_delay_hc_9 : std_logic;
signal measured_delay_hc_7 : std_logic;
signal measured_delay_hc_2 : std_logic;
signal measured_delay_hc_8 : std_logic;
signal measured_delay_hc_12 : std_logic;
signal measured_delay_hc_10 : std_logic;
signal measured_delay_hc_31 : std_logic;
signal measured_delay_hc_11 : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1Z0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_3\ : std_logic;
signal \bfn_8_26_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_11\ : std_logic;
signal \bfn_8_27_0_\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_19\ : std_logic;
signal \bfn_8_28_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \bfn_8_29_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_9_17_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\ : std_logic;
signal \bfn_9_18_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\ : std_logic;
signal \phase_controller_slave.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.N_21\ : std_logic;
signal s3_phy_c : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed11\ : std_logic;
signal \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\ : std_logic;
signal measured_delay_hc_30 : std_logic;
signal measured_delay_hc_24 : std_logic;
signal measured_delay_hc_25 : std_logic;
signal measured_delay_hc_28 : std_logic;
signal measured_delay_hc_29 : std_logic;
signal \delay_measurement_inst.delay_hc_reg3\ : std_logic;
signal measured_delay_hc_23 : std_logic;
signal measured_delay_hc_27 : std_logic;
signal \delay_measurement_inst.un1_elapsed_time_hc\ : std_logic;
signal \delay_measurement_inst.delay_hc_reg3lto31_0_0\ : std_logic;
signal measured_delay_hc_26 : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.elapsed_time_hc_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_136_i_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \bfn_9_26_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_9_27_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_9_28_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_9_29_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_138_i\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \il_max_comp1_D1\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \il_min_comp1_D1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\ : std_logic;
signal measured_delay_tr_15 : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\ : std_logic;
signal \phase_controller_slave.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\ : std_logic;
signal \phase_controller_inst1.stoper_tr.time_passed11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_slave.start_timer_tr_0_sqmuxa\ : std_logic;
signal \il_min_comp2_D1\ : std_logic;
signal \phase_controller_slave.N_20\ : std_logic;
signal \il_min_comp1_D2\ : std_logic;
signal \phase_controller_inst1.T01_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.N_83\ : std_logic;
signal \il_max_comp1_D2\ : std_logic;
signal \phase_controller_inst1.start_timer_hc_0_sqmuxa\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_slave.tr_time_passed\ : std_logic;
signal \phase_controller_slave.stateZ0Z_0\ : std_logic;
signal shift_flag_start : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.N_88\ : std_logic;
signal \il_max_comp2_D2\ : std_logic;
signal \phase_controller_slave.stateZ0Z_4\ : std_logic;
signal \phase_controller_slave.un1_startZ0\ : std_logic;
signal \phase_controller_slave.stateZ0Z_3\ : std_logic;
signal \il_min_comp2_D2\ : std_logic;
signal \phase_controller_slave.stateZ0Z_2\ : std_logic;
signal \phase_controller_slave.hc_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal s2_phy_c : std_logic;
signal \phase_controller_slave.stateZ0Z_1\ : std_logic;
signal s4_phy_c : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.elapsed_time_tr_31\ : std_logic;
signal \delay_measurement_inst.un1_tr_state_1_i_0_0\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.N_86\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_137_i_g\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_3\ : std_logic;
signal s1_phy_c : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_139_i\ : std_logic;
signal delay_tr_input_c : std_logic;
signal delay_tr_d1 : std_logic;
signal delay_tr_d2 : std_logic;
signal \delay_measurement_inst.prev_tr_sigZ0\ : std_logic;
signal \delay_measurement_inst.tr_stateZ0Z_0\ : std_logic;
signal red_c_i : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal delay_hc_input_c : std_logic;
signal delay_hc_d1 : std_logic;
signal \delay_measurement_inst.prev_hc_sigZ0\ : std_logic;
signal \delay_measurement_inst.hc_stateZ0Z_0\ : std_logic;
signal red_c_g : std_logic;
signal delay_hc_d2 : std_logic;
signal clk_100mhz : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_136_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_r_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    reset_wire <= reset;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    il_min_comp1_wire <= il_min_comp1;
    s2_phy <= s2_phy_wire;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_r <= rgb_r_wire;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__12626\,
            RESETB => \N__21350\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__22542\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22544\,
            DIN => \N__22543\,
            DOUT => \N__22542\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22544\,
            PADOUT => \N__22543\,
            PADIN => \N__22542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22533\,
            DIN => \N__22532\,
            DOUT => \N__22531\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22533\,
            PADOUT => \N__22532\,
            PADIN => \N__22531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22524\,
            DIN => \N__22523\,
            DOUT => \N__22522\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22524\,
            PADOUT => \N__22523\,
            PADIN => \N__22522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21530\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22515\,
            DIN => \N__22514\,
            DOUT => \N__22513\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22515\,
            PADOUT => \N__22514\,
            PADIN => \N__22513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21092\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22506\,
            DIN => \N__22505\,
            DOUT => \N__22504\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22506\,
            PADOUT => \N__22505\,
            PADIN => \N__22504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22497\,
            DIN => \N__22496\,
            DOUT => \N__22495\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22497\,
            PADOUT => \N__22496\,
            PADIN => \N__22495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22488\,
            DIN => \N__22487\,
            DOUT => \N__22486\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22488\,
            PADOUT => \N__22487\,
            PADIN => \N__22486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22479\,
            DIN => \N__22478\,
            DOUT => \N__22477\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22479\,
            PADOUT => \N__22478\,
            PADIN => \N__22477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22470\,
            DIN => \N__22469\,
            DOUT => \N__22468\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22470\,
            PADOUT => \N__22469\,
            PADIN => \N__22468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22461\,
            DIN => \N__22460\,
            DOUT => \N__22459\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22461\,
            PADOUT => \N__22460\,
            PADIN => \N__22459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21149\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22452\,
            DIN => \N__22451\,
            DOUT => \N__22450\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__22452\,
            PADOUT => \N__22451\,
            PADIN => \N__22450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18119\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22443\,
            DIN => \N__22442\,
            DOUT => \N__22441\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22443\,
            PADOUT => \N__22442\,
            PADIN => \N__22441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__22434\,
            DIN => \N__22433\,
            DOUT => \N__22432\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__22434\,
            PADOUT => \N__22433\,
            PADIN => \N__22432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5331\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22411\
        );

    \I__5330\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22408\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__22411\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22408\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__5327\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__5325\ : Span12Mux_h
    port map (
            O => \N__22397\,
            I => \N__22394\
        );

    \I__5324\ : Span12Mux_v
    port map (
            O => \N__22394\,
            I => \N__22391\
        );

    \I__5323\ : Odrv12
    port map (
            O => \N__22391\,
            I => delay_hc_input_c
        );

    \I__5322\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22385\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__5320\ : Odrv12
    port map (
            O => \N__22382\,
            I => delay_hc_d1
        );

    \I__5319\ : InMux
    port map (
            O => \N__22379\,
            I => \N__22374\
        );

    \I__5318\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22371\
        );

    \I__5317\ : InMux
    port map (
            O => \N__22377\,
            I => \N__22368\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__22374\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__22371\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__22368\,
            I => \delay_measurement_inst.prev_hc_sigZ0\
        );

    \I__5313\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22356\
        );

    \I__5312\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22353\
        );

    \I__5311\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22350\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__22356\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__22353\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__22350\,
            I => \delay_measurement_inst.hc_stateZ0Z_0\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__22343\,
            I => \N__22336\
        );

    \I__5306\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22332\
        );

    \I__5305\ : InMux
    port map (
            O => \N__22341\,
            I => \N__22329\
        );

    \I__5304\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22326\
        );

    \I__5303\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22323\
        );

    \I__5302\ : InMux
    port map (
            O => \N__22336\,
            I => \N__22320\
        );

    \I__5301\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22317\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__22332\,
            I => \N__22314\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22311\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22308\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22305\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__22320\,
            I => \N__22266\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__22317\,
            I => \N__22244\
        );

    \I__5294\ : Glb2LocalMux
    port map (
            O => \N__22314\,
            I => \N__22082\
        );

    \I__5293\ : Glb2LocalMux
    port map (
            O => \N__22311\,
            I => \N__22082\
        );

    \I__5292\ : Glb2LocalMux
    port map (
            O => \N__22308\,
            I => \N__22082\
        );

    \I__5291\ : Glb2LocalMux
    port map (
            O => \N__22305\,
            I => \N__22082\
        );

    \I__5290\ : SRMux
    port map (
            O => \N__22304\,
            I => \N__22082\
        );

    \I__5289\ : SRMux
    port map (
            O => \N__22303\,
            I => \N__22082\
        );

    \I__5288\ : SRMux
    port map (
            O => \N__22302\,
            I => \N__22082\
        );

    \I__5287\ : SRMux
    port map (
            O => \N__22301\,
            I => \N__22082\
        );

    \I__5286\ : SRMux
    port map (
            O => \N__22300\,
            I => \N__22082\
        );

    \I__5285\ : SRMux
    port map (
            O => \N__22299\,
            I => \N__22082\
        );

    \I__5284\ : SRMux
    port map (
            O => \N__22298\,
            I => \N__22082\
        );

    \I__5283\ : SRMux
    port map (
            O => \N__22297\,
            I => \N__22082\
        );

    \I__5282\ : SRMux
    port map (
            O => \N__22296\,
            I => \N__22082\
        );

    \I__5281\ : SRMux
    port map (
            O => \N__22295\,
            I => \N__22082\
        );

    \I__5280\ : SRMux
    port map (
            O => \N__22294\,
            I => \N__22082\
        );

    \I__5279\ : SRMux
    port map (
            O => \N__22293\,
            I => \N__22082\
        );

    \I__5278\ : SRMux
    port map (
            O => \N__22292\,
            I => \N__22082\
        );

    \I__5277\ : SRMux
    port map (
            O => \N__22291\,
            I => \N__22082\
        );

    \I__5276\ : SRMux
    port map (
            O => \N__22290\,
            I => \N__22082\
        );

    \I__5275\ : SRMux
    port map (
            O => \N__22289\,
            I => \N__22082\
        );

    \I__5274\ : SRMux
    port map (
            O => \N__22288\,
            I => \N__22082\
        );

    \I__5273\ : SRMux
    port map (
            O => \N__22287\,
            I => \N__22082\
        );

    \I__5272\ : SRMux
    port map (
            O => \N__22286\,
            I => \N__22082\
        );

    \I__5271\ : SRMux
    port map (
            O => \N__22285\,
            I => \N__22082\
        );

    \I__5270\ : SRMux
    port map (
            O => \N__22284\,
            I => \N__22082\
        );

    \I__5269\ : SRMux
    port map (
            O => \N__22283\,
            I => \N__22082\
        );

    \I__5268\ : SRMux
    port map (
            O => \N__22282\,
            I => \N__22082\
        );

    \I__5267\ : SRMux
    port map (
            O => \N__22281\,
            I => \N__22082\
        );

    \I__5266\ : SRMux
    port map (
            O => \N__22280\,
            I => \N__22082\
        );

    \I__5265\ : SRMux
    port map (
            O => \N__22279\,
            I => \N__22082\
        );

    \I__5264\ : SRMux
    port map (
            O => \N__22278\,
            I => \N__22082\
        );

    \I__5263\ : SRMux
    port map (
            O => \N__22277\,
            I => \N__22082\
        );

    \I__5262\ : SRMux
    port map (
            O => \N__22276\,
            I => \N__22082\
        );

    \I__5261\ : SRMux
    port map (
            O => \N__22275\,
            I => \N__22082\
        );

    \I__5260\ : SRMux
    port map (
            O => \N__22274\,
            I => \N__22082\
        );

    \I__5259\ : SRMux
    port map (
            O => \N__22273\,
            I => \N__22082\
        );

    \I__5258\ : SRMux
    port map (
            O => \N__22272\,
            I => \N__22082\
        );

    \I__5257\ : SRMux
    port map (
            O => \N__22271\,
            I => \N__22082\
        );

    \I__5256\ : SRMux
    port map (
            O => \N__22270\,
            I => \N__22082\
        );

    \I__5255\ : SRMux
    port map (
            O => \N__22269\,
            I => \N__22082\
        );

    \I__5254\ : Glb2LocalMux
    port map (
            O => \N__22266\,
            I => \N__22082\
        );

    \I__5253\ : SRMux
    port map (
            O => \N__22265\,
            I => \N__22082\
        );

    \I__5252\ : SRMux
    port map (
            O => \N__22264\,
            I => \N__22082\
        );

    \I__5251\ : SRMux
    port map (
            O => \N__22263\,
            I => \N__22082\
        );

    \I__5250\ : SRMux
    port map (
            O => \N__22262\,
            I => \N__22082\
        );

    \I__5249\ : SRMux
    port map (
            O => \N__22261\,
            I => \N__22082\
        );

    \I__5248\ : SRMux
    port map (
            O => \N__22260\,
            I => \N__22082\
        );

    \I__5247\ : SRMux
    port map (
            O => \N__22259\,
            I => \N__22082\
        );

    \I__5246\ : SRMux
    port map (
            O => \N__22258\,
            I => \N__22082\
        );

    \I__5245\ : SRMux
    port map (
            O => \N__22257\,
            I => \N__22082\
        );

    \I__5244\ : SRMux
    port map (
            O => \N__22256\,
            I => \N__22082\
        );

    \I__5243\ : SRMux
    port map (
            O => \N__22255\,
            I => \N__22082\
        );

    \I__5242\ : SRMux
    port map (
            O => \N__22254\,
            I => \N__22082\
        );

    \I__5241\ : SRMux
    port map (
            O => \N__22253\,
            I => \N__22082\
        );

    \I__5240\ : SRMux
    port map (
            O => \N__22252\,
            I => \N__22082\
        );

    \I__5239\ : SRMux
    port map (
            O => \N__22251\,
            I => \N__22082\
        );

    \I__5238\ : SRMux
    port map (
            O => \N__22250\,
            I => \N__22082\
        );

    \I__5237\ : SRMux
    port map (
            O => \N__22249\,
            I => \N__22082\
        );

    \I__5236\ : SRMux
    port map (
            O => \N__22248\,
            I => \N__22082\
        );

    \I__5235\ : SRMux
    port map (
            O => \N__22247\,
            I => \N__22082\
        );

    \I__5234\ : Glb2LocalMux
    port map (
            O => \N__22244\,
            I => \N__22082\
        );

    \I__5233\ : SRMux
    port map (
            O => \N__22243\,
            I => \N__22082\
        );

    \I__5232\ : SRMux
    port map (
            O => \N__22242\,
            I => \N__22082\
        );

    \I__5231\ : SRMux
    port map (
            O => \N__22241\,
            I => \N__22082\
        );

    \I__5230\ : SRMux
    port map (
            O => \N__22240\,
            I => \N__22082\
        );

    \I__5229\ : SRMux
    port map (
            O => \N__22239\,
            I => \N__22082\
        );

    \I__5228\ : SRMux
    port map (
            O => \N__22238\,
            I => \N__22082\
        );

    \I__5227\ : SRMux
    port map (
            O => \N__22237\,
            I => \N__22082\
        );

    \I__5226\ : SRMux
    port map (
            O => \N__22236\,
            I => \N__22082\
        );

    \I__5225\ : SRMux
    port map (
            O => \N__22235\,
            I => \N__22082\
        );

    \I__5224\ : SRMux
    port map (
            O => \N__22234\,
            I => \N__22082\
        );

    \I__5223\ : SRMux
    port map (
            O => \N__22233\,
            I => \N__22082\
        );

    \I__5222\ : SRMux
    port map (
            O => \N__22232\,
            I => \N__22082\
        );

    \I__5221\ : SRMux
    port map (
            O => \N__22231\,
            I => \N__22082\
        );

    \I__5220\ : GlobalMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__5219\ : gio2CtrlBuf
    port map (
            O => \N__22079\,
            I => red_c_g
        );

    \I__5218\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22072\
        );

    \I__5217\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22067\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__22072\,
            I => \N__22064\
        );

    \I__5215\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22061\
        );

    \I__5214\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22058\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22051\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__22064\,
            I => \N__22051\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22051\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22048\
        );

    \I__5209\ : Odrv4
    port map (
            O => \N__22051\,
            I => delay_hc_d2
        );

    \I__5208\ : Odrv12
    port map (
            O => \N__22048\,
            I => delay_hc_d2
        );

    \I__5207\ : ClkMux
    port map (
            O => \N__22043\,
            I => \N__21788\
        );

    \I__5206\ : ClkMux
    port map (
            O => \N__22042\,
            I => \N__21788\
        );

    \I__5205\ : ClkMux
    port map (
            O => \N__22041\,
            I => \N__21788\
        );

    \I__5204\ : ClkMux
    port map (
            O => \N__22040\,
            I => \N__21788\
        );

    \I__5203\ : ClkMux
    port map (
            O => \N__22039\,
            I => \N__21788\
        );

    \I__5202\ : ClkMux
    port map (
            O => \N__22038\,
            I => \N__21788\
        );

    \I__5201\ : ClkMux
    port map (
            O => \N__22037\,
            I => \N__21788\
        );

    \I__5200\ : ClkMux
    port map (
            O => \N__22036\,
            I => \N__21788\
        );

    \I__5199\ : ClkMux
    port map (
            O => \N__22035\,
            I => \N__21788\
        );

    \I__5198\ : ClkMux
    port map (
            O => \N__22034\,
            I => \N__21788\
        );

    \I__5197\ : ClkMux
    port map (
            O => \N__22033\,
            I => \N__21788\
        );

    \I__5196\ : ClkMux
    port map (
            O => \N__22032\,
            I => \N__21788\
        );

    \I__5195\ : ClkMux
    port map (
            O => \N__22031\,
            I => \N__21788\
        );

    \I__5194\ : ClkMux
    port map (
            O => \N__22030\,
            I => \N__21788\
        );

    \I__5193\ : ClkMux
    port map (
            O => \N__22029\,
            I => \N__21788\
        );

    \I__5192\ : ClkMux
    port map (
            O => \N__22028\,
            I => \N__21788\
        );

    \I__5191\ : ClkMux
    port map (
            O => \N__22027\,
            I => \N__21788\
        );

    \I__5190\ : ClkMux
    port map (
            O => \N__22026\,
            I => \N__21788\
        );

    \I__5189\ : ClkMux
    port map (
            O => \N__22025\,
            I => \N__21788\
        );

    \I__5188\ : ClkMux
    port map (
            O => \N__22024\,
            I => \N__21788\
        );

    \I__5187\ : ClkMux
    port map (
            O => \N__22023\,
            I => \N__21788\
        );

    \I__5186\ : ClkMux
    port map (
            O => \N__22022\,
            I => \N__21788\
        );

    \I__5185\ : ClkMux
    port map (
            O => \N__22021\,
            I => \N__21788\
        );

    \I__5184\ : ClkMux
    port map (
            O => \N__22020\,
            I => \N__21788\
        );

    \I__5183\ : ClkMux
    port map (
            O => \N__22019\,
            I => \N__21788\
        );

    \I__5182\ : ClkMux
    port map (
            O => \N__22018\,
            I => \N__21788\
        );

    \I__5181\ : ClkMux
    port map (
            O => \N__22017\,
            I => \N__21788\
        );

    \I__5180\ : ClkMux
    port map (
            O => \N__22016\,
            I => \N__21788\
        );

    \I__5179\ : ClkMux
    port map (
            O => \N__22015\,
            I => \N__21788\
        );

    \I__5178\ : ClkMux
    port map (
            O => \N__22014\,
            I => \N__21788\
        );

    \I__5177\ : ClkMux
    port map (
            O => \N__22013\,
            I => \N__21788\
        );

    \I__5176\ : ClkMux
    port map (
            O => \N__22012\,
            I => \N__21788\
        );

    \I__5175\ : ClkMux
    port map (
            O => \N__22011\,
            I => \N__21788\
        );

    \I__5174\ : ClkMux
    port map (
            O => \N__22010\,
            I => \N__21788\
        );

    \I__5173\ : ClkMux
    port map (
            O => \N__22009\,
            I => \N__21788\
        );

    \I__5172\ : ClkMux
    port map (
            O => \N__22008\,
            I => \N__21788\
        );

    \I__5171\ : ClkMux
    port map (
            O => \N__22007\,
            I => \N__21788\
        );

    \I__5170\ : ClkMux
    port map (
            O => \N__22006\,
            I => \N__21788\
        );

    \I__5169\ : ClkMux
    port map (
            O => \N__22005\,
            I => \N__21788\
        );

    \I__5168\ : ClkMux
    port map (
            O => \N__22004\,
            I => \N__21788\
        );

    \I__5167\ : ClkMux
    port map (
            O => \N__22003\,
            I => \N__21788\
        );

    \I__5166\ : ClkMux
    port map (
            O => \N__22002\,
            I => \N__21788\
        );

    \I__5165\ : ClkMux
    port map (
            O => \N__22001\,
            I => \N__21788\
        );

    \I__5164\ : ClkMux
    port map (
            O => \N__22000\,
            I => \N__21788\
        );

    \I__5163\ : ClkMux
    port map (
            O => \N__21999\,
            I => \N__21788\
        );

    \I__5162\ : ClkMux
    port map (
            O => \N__21998\,
            I => \N__21788\
        );

    \I__5161\ : ClkMux
    port map (
            O => \N__21997\,
            I => \N__21788\
        );

    \I__5160\ : ClkMux
    port map (
            O => \N__21996\,
            I => \N__21788\
        );

    \I__5159\ : ClkMux
    port map (
            O => \N__21995\,
            I => \N__21788\
        );

    \I__5158\ : ClkMux
    port map (
            O => \N__21994\,
            I => \N__21788\
        );

    \I__5157\ : ClkMux
    port map (
            O => \N__21993\,
            I => \N__21788\
        );

    \I__5156\ : ClkMux
    port map (
            O => \N__21992\,
            I => \N__21788\
        );

    \I__5155\ : ClkMux
    port map (
            O => \N__21991\,
            I => \N__21788\
        );

    \I__5154\ : ClkMux
    port map (
            O => \N__21990\,
            I => \N__21788\
        );

    \I__5153\ : ClkMux
    port map (
            O => \N__21989\,
            I => \N__21788\
        );

    \I__5152\ : ClkMux
    port map (
            O => \N__21988\,
            I => \N__21788\
        );

    \I__5151\ : ClkMux
    port map (
            O => \N__21987\,
            I => \N__21788\
        );

    \I__5150\ : ClkMux
    port map (
            O => \N__21986\,
            I => \N__21788\
        );

    \I__5149\ : ClkMux
    port map (
            O => \N__21985\,
            I => \N__21788\
        );

    \I__5148\ : ClkMux
    port map (
            O => \N__21984\,
            I => \N__21788\
        );

    \I__5147\ : ClkMux
    port map (
            O => \N__21983\,
            I => \N__21788\
        );

    \I__5146\ : ClkMux
    port map (
            O => \N__21982\,
            I => \N__21788\
        );

    \I__5145\ : ClkMux
    port map (
            O => \N__21981\,
            I => \N__21788\
        );

    \I__5144\ : ClkMux
    port map (
            O => \N__21980\,
            I => \N__21788\
        );

    \I__5143\ : ClkMux
    port map (
            O => \N__21979\,
            I => \N__21788\
        );

    \I__5142\ : ClkMux
    port map (
            O => \N__21978\,
            I => \N__21788\
        );

    \I__5141\ : ClkMux
    port map (
            O => \N__21977\,
            I => \N__21788\
        );

    \I__5140\ : ClkMux
    port map (
            O => \N__21976\,
            I => \N__21788\
        );

    \I__5139\ : ClkMux
    port map (
            O => \N__21975\,
            I => \N__21788\
        );

    \I__5138\ : ClkMux
    port map (
            O => \N__21974\,
            I => \N__21788\
        );

    \I__5137\ : ClkMux
    port map (
            O => \N__21973\,
            I => \N__21788\
        );

    \I__5136\ : ClkMux
    port map (
            O => \N__21972\,
            I => \N__21788\
        );

    \I__5135\ : ClkMux
    port map (
            O => \N__21971\,
            I => \N__21788\
        );

    \I__5134\ : ClkMux
    port map (
            O => \N__21970\,
            I => \N__21788\
        );

    \I__5133\ : ClkMux
    port map (
            O => \N__21969\,
            I => \N__21788\
        );

    \I__5132\ : ClkMux
    port map (
            O => \N__21968\,
            I => \N__21788\
        );

    \I__5131\ : ClkMux
    port map (
            O => \N__21967\,
            I => \N__21788\
        );

    \I__5130\ : ClkMux
    port map (
            O => \N__21966\,
            I => \N__21788\
        );

    \I__5129\ : ClkMux
    port map (
            O => \N__21965\,
            I => \N__21788\
        );

    \I__5128\ : ClkMux
    port map (
            O => \N__21964\,
            I => \N__21788\
        );

    \I__5127\ : ClkMux
    port map (
            O => \N__21963\,
            I => \N__21788\
        );

    \I__5126\ : ClkMux
    port map (
            O => \N__21962\,
            I => \N__21788\
        );

    \I__5125\ : ClkMux
    port map (
            O => \N__21961\,
            I => \N__21788\
        );

    \I__5124\ : ClkMux
    port map (
            O => \N__21960\,
            I => \N__21788\
        );

    \I__5123\ : ClkMux
    port map (
            O => \N__21959\,
            I => \N__21788\
        );

    \I__5122\ : GlobalMux
    port map (
            O => \N__21788\,
            I => clk_100mhz
        );

    \I__5121\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__21782\,
            I => \N__21778\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21781\,
            I => \N__21774\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__21778\,
            I => \N__21771\
        );

    \I__5117\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21768\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__21774\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__21771\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__21768\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21761\,
            I => \N__21756\
        );

    \I__5112\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21752\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21749\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__21756\,
            I => \N__21746\
        );

    \I__5109\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21743\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__21752\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__21749\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__21746\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__21743\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__5104\ : IoInMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__5102\ : Odrv12
    port map (
            O => \N__21728\,
            I => \delay_measurement_inst.delay_hc_timer.N_136_i\
        );

    \I__5101\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21722\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21722\,
            I => \N__21718\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21715\
        );

    \I__5098\ : Span4Mux_s1_v
    port map (
            O => \N__21718\,
            I => \N__21710\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21710\
        );

    \I__5096\ : Span4Mux_v
    port map (
            O => \N__21710\,
            I => \N__21704\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21701\
        );

    \I__5094\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21698\
        );

    \I__5093\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21695\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__21704\,
            I => \N__21692\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21687\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__21698\,
            I => \N__21687\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21695\,
            I => \N__21684\
        );

    \I__5088\ : Sp12to4
    port map (
            O => \N__21692\,
            I => \N__21681\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__21687\,
            I => \N__21678\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__21684\,
            I => \N__21675\
        );

    \I__5085\ : Span12Mux_v
    port map (
            O => \N__21681\,
            I => \N__21672\
        );

    \I__5084\ : Sp12to4
    port map (
            O => \N__21678\,
            I => \N__21669\
        );

    \I__5083\ : Span4Mux_h
    port map (
            O => \N__21675\,
            I => \N__21666\
        );

    \I__5082\ : Span12Mux_v
    port map (
            O => \N__21672\,
            I => \N__21663\
        );

    \I__5081\ : Span12Mux_h
    port map (
            O => \N__21669\,
            I => \N__21660\
        );

    \I__5080\ : Sp12to4
    port map (
            O => \N__21666\,
            I => \N__21657\
        );

    \I__5079\ : Span12Mux_h
    port map (
            O => \N__21663\,
            I => \N__21652\
        );

    \I__5078\ : Span12Mux_v
    port map (
            O => \N__21660\,
            I => \N__21652\
        );

    \I__5077\ : Span12Mux_v
    port map (
            O => \N__21657\,
            I => \N__21649\
        );

    \I__5076\ : Odrv12
    port map (
            O => \N__21652\,
            I => start_stop_c
        );

    \I__5075\ : Odrv12
    port map (
            O => \N__21649\,
            I => start_stop_c
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__21644\,
            I => \N__21639\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21630\
        );

    \I__5072\ : InMux
    port map (
            O => \N__21642\,
            I => \N__21630\
        );

    \I__5071\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21630\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21627\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21624\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__21630\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__21627\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__21624\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__21611\,
            I => \phase_controller_inst1.N_86\
        );

    \I__5062\ : CEMux
    port map (
            O => \N__21608\,
            I => \N__21603\
        );

    \I__5061\ : CEMux
    port map (
            O => \N__21607\,
            I => \N__21600\
        );

    \I__5060\ : CEMux
    port map (
            O => \N__21606\,
            I => \N__21597\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21603\,
            I => \N__21593\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__21600\,
            I => \N__21590\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__21597\,
            I => \N__21587\
        );

    \I__5056\ : CEMux
    port map (
            O => \N__21596\,
            I => \N__21584\
        );

    \I__5055\ : Span4Mux_h
    port map (
            O => \N__21593\,
            I => \N__21581\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__21590\,
            I => \N__21578\
        );

    \I__5053\ : Span4Mux_h
    port map (
            O => \N__21587\,
            I => \N__21575\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__21584\,
            I => \N__21572\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__21581\,
            I => \delay_measurement_inst.delay_hc_timer.N_137_i_g\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__21578\,
            I => \delay_measurement_inst.delay_hc_timer.N_137_i_g\
        );

    \I__5049\ : Odrv4
    port map (
            O => \N__21575\,
            I => \delay_measurement_inst.delay_hc_timer.N_137_i_g\
        );

    \I__5048\ : Odrv12
    port map (
            O => \N__21572\,
            I => \delay_measurement_inst.delay_hc_timer.N_137_i_g\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21563\,
            I => \N__21560\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__5045\ : Span4Mux_v
    port map (
            O => \N__21557\,
            I => \N__21553\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__21556\,
            I => \N__21549\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__21553\,
            I => \N__21545\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21552\,
            I => \N__21540\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21540\
        );

    \I__5040\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21537\
        );

    \I__5039\ : Odrv4
    port map (
            O => \N__21545\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21540\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__21537\,
            I => \phase_controller_inst1.stateZ0Z_3\
        );

    \I__5036\ : IoInMux
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__5034\ : Span4Mux_s3_v
    port map (
            O => \N__21524\,
            I => \N__21521\
        );

    \I__5033\ : Span4Mux_h
    port map (
            O => \N__21521\,
            I => \N__21518\
        );

    \I__5032\ : Odrv4
    port map (
            O => \N__21518\,
            I => s1_phy_c
        );

    \I__5031\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21510\
        );

    \I__5030\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21507\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21504\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21510\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21507\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__21504\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21493\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21490\
        );

    \I__5023\ : LocalMux
    port map (
            O => \N__21493\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21490\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__5021\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21481\
        );

    \I__5020\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21476\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21473\
        );

    \I__5018\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21470\
        );

    \I__5017\ : InMux
    port map (
            O => \N__21479\,
            I => \N__21467\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__21476\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5015\ : Odrv12
    port map (
            O => \N__21473\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21470\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5013\ : LocalMux
    port map (
            O => \N__21467\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__5012\ : IoInMux
    port map (
            O => \N__21458\,
            I => \N__21455\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__21455\,
            I => \N__21452\
        );

    \I__5010\ : Span12Mux_s2_v
    port map (
            O => \N__21452\,
            I => \N__21449\
        );

    \I__5009\ : Odrv12
    port map (
            O => \N__21449\,
            I => \delay_measurement_inst.delay_tr_timer.N_139_i\
        );

    \I__5008\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21443\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21440\
        );

    \I__5006\ : Span4Mux_h
    port map (
            O => \N__21440\,
            I => \N__21437\
        );

    \I__5005\ : Span4Mux_v
    port map (
            O => \N__21437\,
            I => \N__21434\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__21434\,
            I => \N__21431\
        );

    \I__5003\ : Odrv4
    port map (
            O => \N__21431\,
            I => delay_tr_input_c
        );

    \I__5002\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21425\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__21425\,
            I => delay_tr_d1
        );

    \I__5000\ : CascadeMux
    port map (
            O => \N__21422\,
            I => \N__21415\
        );

    \I__4999\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21412\
        );

    \I__4998\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21405\
        );

    \I__4997\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21405\
        );

    \I__4996\ : InMux
    port map (
            O => \N__21418\,
            I => \N__21405\
        );

    \I__4995\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21402\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__21412\,
            I => delay_tr_d2
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__21405\,
            I => delay_tr_d2
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__21402\,
            I => delay_tr_d2
        );

    \I__4991\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21389\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21384\
        );

    \I__4989\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21384\
        );

    \I__4988\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21381\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21389\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21384\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__21381\,
            I => \delay_measurement_inst.prev_tr_sigZ0\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__4983\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21365\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21362\
        );

    \I__4981\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21359\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__21368\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__21365\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__21362\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__21359\,
            I => \delay_measurement_inst.tr_stateZ0Z_0\
        );

    \I__4976\ : IoInMux
    port map (
            O => \N__21350\,
            I => \N__21346\
        );

    \I__4975\ : CEMux
    port map (
            O => \N__21349\,
            I => \N__21343\
        );

    \I__4974\ : LocalMux
    port map (
            O => \N__21346\,
            I => \N__21339\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21343\,
            I => \N__21335\
        );

    \I__4972\ : CEMux
    port map (
            O => \N__21342\,
            I => \N__21332\
        );

    \I__4971\ : IoSpan4Mux
    port map (
            O => \N__21339\,
            I => \N__21328\
        );

    \I__4970\ : CEMux
    port map (
            O => \N__21338\,
            I => \N__21325\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__21335\,
            I => \N__21319\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21319\
        );

    \I__4967\ : CEMux
    port map (
            O => \N__21331\,
            I => \N__21316\
        );

    \I__4966\ : Span4Mux_s2_v
    port map (
            O => \N__21328\,
            I => \N__21312\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__21325\,
            I => \N__21309\
        );

    \I__4964\ : CEMux
    port map (
            O => \N__21324\,
            I => \N__21306\
        );

    \I__4963\ : Span4Mux_v
    port map (
            O => \N__21319\,
            I => \N__21301\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21301\
        );

    \I__4961\ : CEMux
    port map (
            O => \N__21315\,
            I => \N__21298\
        );

    \I__4960\ : Span4Mux_h
    port map (
            O => \N__21312\,
            I => \N__21293\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__21309\,
            I => \N__21293\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__21306\,
            I => \N__21290\
        );

    \I__4957\ : Span4Mux_h
    port map (
            O => \N__21301\,
            I => \N__21286\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21283\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__21293\,
            I => \N__21278\
        );

    \I__4954\ : Span4Mux_v
    port map (
            O => \N__21290\,
            I => \N__21278\
        );

    \I__4953\ : CEMux
    port map (
            O => \N__21289\,
            I => \N__21275\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__21286\,
            I => \N__21270\
        );

    \I__4951\ : Span4Mux_v
    port map (
            O => \N__21283\,
            I => \N__21270\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__21278\,
            I => \N__21267\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__21275\,
            I => \N__21264\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__21270\,
            I => \N__21261\
        );

    \I__4947\ : Span4Mux_h
    port map (
            O => \N__21267\,
            I => \N__21258\
        );

    \I__4946\ : Span4Mux_v
    port map (
            O => \N__21264\,
            I => \N__21255\
        );

    \I__4945\ : Odrv4
    port map (
            O => \N__21261\,
            I => red_c_i
        );

    \I__4944\ : Odrv4
    port map (
            O => \N__21258\,
            I => red_c_i
        );

    \I__4943\ : Odrv4
    port map (
            O => \N__21255\,
            I => red_c_i
        );

    \I__4942\ : InMux
    port map (
            O => \N__21248\,
            I => \N__21244\
        );

    \I__4941\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__21244\,
            I => \N__21235\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__21241\,
            I => \N__21235\
        );

    \I__4938\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21232\
        );

    \I__4937\ : Odrv12
    port map (
            O => \N__21235\,
            I => \il_min_comp2_D2\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__21232\,
            I => \il_min_comp2_D2\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__21227\,
            I => \N__21223\
        );

    \I__4934\ : InMux
    port map (
            O => \N__21226\,
            I => \N__21219\
        );

    \I__4933\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21216\
        );

    \I__4932\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21213\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__21219\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__21216\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__21213\,
            I => \phase_controller_slave.stateZ0Z_2\
        );

    \I__4928\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21200\
        );

    \I__4927\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21197\
        );

    \I__4926\ : InMux
    port map (
            O => \N__21204\,
            I => \N__21194\
        );

    \I__4925\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21191\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__21200\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__21197\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__21194\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__21191\,
            I => \phase_controller_slave.hc_time_passed\
        );

    \I__4920\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21177\
        );

    \I__4919\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21174\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__21180\,
            I => \N__21171\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__21177\,
            I => \N__21167\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21164\
        );

    \I__4915\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21161\
        );

    \I__4914\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21158\
        );

    \I__4913\ : Odrv12
    port map (
            O => \N__21167\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__21164\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__21161\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__21158\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__4909\ : IoInMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__4907\ : Span4Mux_s0_v
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__4906\ : Span4Mux_v
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__4905\ : Span4Mux_v
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__21134\,
            I => s2_phy_c
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__21131\,
            I => \N__21127\
        );

    \I__4902\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21122\
        );

    \I__4901\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21119\
        );

    \I__4900\ : CascadeMux
    port map (
            O => \N__21126\,
            I => \N__21116\
        );

    \I__4899\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21113\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__21122\,
            I => \N__21110\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21107\
        );

    \I__4896\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21104\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N__21101\
        );

    \I__4894\ : Odrv12
    port map (
            O => \N__21110\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__21107\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__21104\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__4891\ : Odrv12
    port map (
            O => \N__21101\,
            I => \phase_controller_slave.stateZ0Z_1\
        );

    \I__4890\ : IoInMux
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__4888\ : Span4Mux_s1_v
    port map (
            O => \N__21086\,
            I => \N__21083\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__21080\,
            I => s4_phy_c
        );

    \I__4885\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21067\
        );

    \I__4884\ : InMux
    port map (
            O => \N__21076\,
            I => \N__21067\
        );

    \I__4883\ : InMux
    port map (
            O => \N__21075\,
            I => \N__21046\
        );

    \I__4882\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21046\
        );

    \I__4881\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21046\
        );

    \I__4880\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21046\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__21067\,
            I => \N__21031\
        );

    \I__4878\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21022\
        );

    \I__4877\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21022\
        );

    \I__4876\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21022\
        );

    \I__4875\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21022\
        );

    \I__4874\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21013\
        );

    \I__4873\ : InMux
    port map (
            O => \N__21061\,
            I => \N__21013\
        );

    \I__4872\ : InMux
    port map (
            O => \N__21060\,
            I => \N__21013\
        );

    \I__4871\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21013\
        );

    \I__4870\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21004\
        );

    \I__4869\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21004\
        );

    \I__4868\ : InMux
    port map (
            O => \N__21056\,
            I => \N__21004\
        );

    \I__4867\ : InMux
    port map (
            O => \N__21055\,
            I => \N__21004\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__21046\,
            I => \N__21001\
        );

    \I__4865\ : InMux
    port map (
            O => \N__21045\,
            I => \N__20992\
        );

    \I__4864\ : InMux
    port map (
            O => \N__21044\,
            I => \N__20992\
        );

    \I__4863\ : InMux
    port map (
            O => \N__21043\,
            I => \N__20992\
        );

    \I__4862\ : InMux
    port map (
            O => \N__21042\,
            I => \N__20992\
        );

    \I__4861\ : InMux
    port map (
            O => \N__21041\,
            I => \N__20983\
        );

    \I__4860\ : InMux
    port map (
            O => \N__21040\,
            I => \N__20983\
        );

    \I__4859\ : InMux
    port map (
            O => \N__21039\,
            I => \N__20983\
        );

    \I__4858\ : InMux
    port map (
            O => \N__21038\,
            I => \N__20983\
        );

    \I__4857\ : InMux
    port map (
            O => \N__21037\,
            I => \N__20974\
        );

    \I__4856\ : InMux
    port map (
            O => \N__21036\,
            I => \N__20974\
        );

    \I__4855\ : InMux
    port map (
            O => \N__21035\,
            I => \N__20974\
        );

    \I__4854\ : InMux
    port map (
            O => \N__21034\,
            I => \N__20974\
        );

    \I__4853\ : Span4Mux_h
    port map (
            O => \N__21031\,
            I => \N__20969\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__21022\,
            I => \N__20969\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__21013\,
            I => \N__20962\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__21004\,
            I => \N__20962\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__21001\,
            I => \N__20962\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__20992\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__20983\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__20974\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4845\ : Odrv4
    port map (
            O => \N__20969\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4844\ : Odrv4
    port map (
            O => \N__20962\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__4843\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20948\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__20948\,
            I => \N__20932\
        );

    \I__4841\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20921\
        );

    \I__4840\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20921\
        );

    \I__4839\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20921\
        );

    \I__4838\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20921\
        );

    \I__4837\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20921\
        );

    \I__4836\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20914\
        );

    \I__4835\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20914\
        );

    \I__4834\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20914\
        );

    \I__4833\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20907\
        );

    \I__4832\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20907\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20937\,
            I => \N__20907\
        );

    \I__4830\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20902\
        );

    \I__4829\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20902\
        );

    \I__4828\ : Span4Mux_h
    port map (
            O => \N__20932\,
            I => \N__20899\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__20921\,
            I => \N__20896\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__20914\,
            I => \N__20889\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__20907\,
            I => \N__20889\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__20902\,
            I => \N__20889\
        );

    \I__4823\ : Span4Mux_v
    port map (
            O => \N__20899\,
            I => \N__20886\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__20896\,
            I => \N__20881\
        );

    \I__4821\ : Span4Mux_v
    port map (
            O => \N__20889\,
            I => \N__20881\
        );

    \I__4820\ : Span4Mux_h
    port map (
            O => \N__20886\,
            I => \N__20878\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__20881\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__20878\,
            I => \delay_measurement_inst.elapsed_time_tr_31\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__4816\ : InMux
    port map (
            O => \N__20870\,
            I => \N__20867\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__20867\,
            I => \N__20864\
        );

    \I__4814\ : Span4Mux_h
    port map (
            O => \N__20864\,
            I => \N__20861\
        );

    \I__4813\ : Span4Mux_h
    port map (
            O => \N__20861\,
            I => \N__20858\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__20858\,
            I => \delay_measurement_inst.un1_tr_state_1_i_0_0\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20849\
        );

    \I__4810\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20849\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__20849\,
            I => \phase_controller_inst1.T01_0_sqmuxa\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__20846\,
            I => \N__20834\
        );

    \I__4807\ : CascadeMux
    port map (
            O => \N__20845\,
            I => \N__20831\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__20844\,
            I => \N__20828\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__20843\,
            I => \N__20821\
        );

    \I__4804\ : CascadeMux
    port map (
            O => \N__20842\,
            I => \N__20818\
        );

    \I__4803\ : CascadeMux
    port map (
            O => \N__20841\,
            I => \N__20815\
        );

    \I__4802\ : CascadeMux
    port map (
            O => \N__20840\,
            I => \N__20805\
        );

    \I__4801\ : CascadeMux
    port map (
            O => \N__20839\,
            I => \N__20802\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__20838\,
            I => \N__20799\
        );

    \I__4799\ : CascadeMux
    port map (
            O => \N__20837\,
            I => \N__20796\
        );

    \I__4798\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20781\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20831\,
            I => \N__20781\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20781\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20827\,
            I => \N__20781\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20826\,
            I => \N__20781\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20781\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20781\
        );

    \I__4791\ : InMux
    port map (
            O => \N__20821\,
            I => \N__20775\
        );

    \I__4790\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20766\
        );

    \I__4789\ : InMux
    port map (
            O => \N__20815\,
            I => \N__20766\
        );

    \I__4788\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20766\
        );

    \I__4787\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20766\
        );

    \I__4786\ : CascadeMux
    port map (
            O => \N__20812\,
            I => \N__20763\
        );

    \I__4785\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20746\
        );

    \I__4784\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20746\
        );

    \I__4783\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20746\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20746\
        );

    \I__4781\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20746\
        );

    \I__4780\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20746\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20746\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20746\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20743\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20738\
        );

    \I__4775\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20738\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__20778\,
            I => \N__20735\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__20775\,
            I => \N__20730\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20766\,
            I => \N__20730\
        );

    \I__4771\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20727\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__20746\,
            I => \N__20724\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__20743\,
            I => \N__20721\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20718\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20735\,
            I => \N__20715\
        );

    \I__4766\ : Span4Mux_v
    port map (
            O => \N__20730\,
            I => \N__20712\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__20727\,
            I => \N__20707\
        );

    \I__4764\ : Span4Mux_h
    port map (
            O => \N__20724\,
            I => \N__20707\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__20721\,
            I => \N__20704\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__20718\,
            I => \N__20701\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20715\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__20712\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__20707\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__20704\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__20701\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__4756\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20684\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20684\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20684\,
            I => \phase_controller_inst1.N_83\
        );

    \I__4753\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20674\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20680\,
            I => \N__20674\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20671\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__20674\,
            I => \N__20666\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__20671\,
            I => \N__20666\
        );

    \I__4748\ : Odrv12
    port map (
            O => \N__20666\,
            I => \il_max_comp1_D2\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__20660\,
            I => \phase_controller_inst1.start_timer_hc_0_sqmuxa\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__20657\,
            I => \N__20641\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__20656\,
            I => \N__20638\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__20655\,
            I => \N__20635\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \N__20629\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__20653\,
            I => \N__20626\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__20652\,
            I => \N__20623\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__20651\,
            I => \N__20620\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \N__20617\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__20649\,
            I => \N__20612\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__20648\,
            I => \N__20608\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__20647\,
            I => \N__20605\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__20646\,
            I => \N__20602\
        );

    \I__4733\ : CascadeMux
    port map (
            O => \N__20645\,
            I => \N__20599\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__20644\,
            I => \N__20596\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20581\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20638\,
            I => \N__20581\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20581\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20581\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20581\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20581\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20572\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20572\
        );

    \I__4723\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20572\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20572\
        );

    \I__4721\ : InMux
    port map (
            O => \N__20617\,
            I => \N__20565\
        );

    \I__4720\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20565\
        );

    \I__4719\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20565\
        );

    \I__4718\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20560\
        );

    \I__4717\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20560\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20551\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20551\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20551\
        );

    \I__4713\ : InMux
    port map (
            O => \N__20599\,
            I => \N__20551\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20546\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20546\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20542\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20539\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__20572\,
            I => \N__20534\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20565\,
            I => \N__20534\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__20560\,
            I => \N__20527\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20527\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__20546\,
            I => \N__20527\
        );

    \I__4703\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20524\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20520\
        );

    \I__4701\ : Span4Mux_h
    port map (
            O => \N__20539\,
            I => \N__20513\
        );

    \I__4700\ : Span4Mux_v
    port map (
            O => \N__20534\,
            I => \N__20513\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__20527\,
            I => \N__20513\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20524\,
            I => \N__20510\
        );

    \I__4697\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20507\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20520\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__20513\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__20510\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__20507\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20491\
        );

    \I__4691\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20496\,
            I => \N__20488\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20491\,
            I => \N__20484\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N__20481\
        );

    \I__4687\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20478\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__20484\,
            I => \N__20475\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__20481\,
            I => \N__20472\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__20478\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__4683\ : Odrv4
    port map (
            O => \N__20475\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__20472\,
            I => \phase_controller_slave.tr_time_passed\
        );

    \I__4681\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20458\
        );

    \I__4680\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20458\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20455\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__20458\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__20455\,
            I => \phase_controller_slave.stateZ0Z_0\
        );

    \I__4676\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20446\
        );

    \I__4675\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__20446\,
            I => shift_flag_start
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__20443\,
            I => shift_flag_start
        );

    \I__4672\ : InMux
    port map (
            O => \N__20438\,
            I => \N__20432\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20437\,
            I => \N__20427\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20436\,
            I => \N__20427\
        );

    \I__4669\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20424\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__20432\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20427\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__20424\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20411\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20411\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20407\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20404\
        );

    \I__4661\ : Span4Mux_h
    port map (
            O => \N__20407\,
            I => \N__20400\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20404\,
            I => \N__20397\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20394\
        );

    \I__4658\ : Sp12to4
    port map (
            O => \N__20400\,
            I => \N__20391\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__20397\,
            I => \N__20388\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__20394\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__4655\ : Odrv12
    port map (
            O => \N__20391\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__20388\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20378\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20378\,
            I => \phase_controller_inst1.N_88\
        );

    \I__4651\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20369\
        );

    \I__4650\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20369\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__20369\,
            I => \N__20366\
        );

    \I__4648\ : Span4Mux_h
    port map (
            O => \N__20366\,
            I => \N__20362\
        );

    \I__4647\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20359\
        );

    \I__4646\ : Sp12to4
    port map (
            O => \N__20362\,
            I => \N__20354\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__20359\,
            I => \N__20354\
        );

    \I__4644\ : Span12Mux_v
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__4643\ : Odrv12
    port map (
            O => \N__20351\,
            I => \il_max_comp2_D2\
        );

    \I__4642\ : CascadeMux
    port map (
            O => \N__20348\,
            I => \N__20345\
        );

    \I__4641\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20340\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__20344\,
            I => \N__20337\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__20343\,
            I => \N__20334\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__20340\,
            I => \N__20330\
        );

    \I__4637\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20327\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20324\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__20333\,
            I => \N__20321\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__20330\,
            I => \N__20318\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20315\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20312\
        );

    \I__4631\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20309\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__20318\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__20315\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__20312\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20309\,
            I => \phase_controller_slave.stateZ0Z_4\
        );

    \I__4626\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20296\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20293\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__20296\,
            I => \phase_controller_slave.un1_startZ0\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__20293\,
            I => \phase_controller_slave.un1_startZ0\
        );

    \I__4622\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20282\
        );

    \I__4621\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20277\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20277\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20285\,
            I => \N__20274\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__20282\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20277\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__20274\,
            I => \phase_controller_slave.stateZ0Z_3\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__20267\,
            I => \N__20263\
        );

    \I__4614\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20257\
        );

    \I__4613\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20257\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20254\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__20257\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__20254\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__4609\ : InMux
    port map (
            O => \N__20249\,
            I => \N__20245\
        );

    \I__4608\ : InMux
    port map (
            O => \N__20248\,
            I => \N__20242\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__20245\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__20242\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__4605\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20234\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__20234\,
            I => \phase_controller_slave.start_timer_tr_0_sqmuxa\
        );

    \I__4603\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__20228\,
            I => \N__20225\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__20225\,
            I => \N__20222\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__4599\ : Odrv4
    port map (
            O => \N__20219\,
            I => \il_min_comp2_D1\
        );

    \I__4598\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20213\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__20213\,
            I => \phase_controller_slave.N_20\
        );

    \I__4596\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20205\
        );

    \I__4595\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20202\
        );

    \I__4594\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20199\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__20205\,
            I => \N__20196\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20191\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__20199\,
            I => \N__20191\
        );

    \I__4590\ : Odrv12
    port map (
            O => \N__20196\,
            I => \il_min_comp1_D2\
        );

    \I__4589\ : Odrv4
    port map (
            O => \N__20191\,
            I => \il_min_comp1_D2\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__4586\ : Span4Mux_h
    port map (
            O => \N__20180\,
            I => \N__20177\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__20177\,
            I => \N__20174\
        );

    \I__4584\ : Span4Mux_v
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__20171\,
            I => il_max_comp1_c
        );

    \I__4582\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20165\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__20165\,
            I => \il_max_comp1_D1\
        );

    \I__4580\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__20159\,
            I => \N__20156\
        );

    \I__4578\ : Span4Mux_v
    port map (
            O => \N__20156\,
            I => \N__20153\
        );

    \I__4577\ : Sp12to4
    port map (
            O => \N__20153\,
            I => \N__20150\
        );

    \I__4576\ : Span12Mux_h
    port map (
            O => \N__20150\,
            I => \N__20147\
        );

    \I__4575\ : Odrv12
    port map (
            O => \N__20147\,
            I => il_min_comp1_c
        );

    \I__4574\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20141\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__20141\,
            I => \il_min_comp1_D1\
        );

    \I__4572\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20132\
        );

    \I__4571\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20121\
        );

    \I__4570\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20121\
        );

    \I__4569\ : InMux
    port map (
            O => \N__20135\,
            I => \N__20121\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__20132\,
            I => \N__20113\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__20131\,
            I => \N__20110\
        );

    \I__4566\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20104\
        );

    \I__4565\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20104\
        );

    \I__4564\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20101\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__20121\,
            I => \N__20098\
        );

    \I__4562\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20089\
        );

    \I__4561\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20089\
        );

    \I__4560\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20089\
        );

    \I__4559\ : InMux
    port map (
            O => \N__20117\,
            I => \N__20089\
        );

    \I__4558\ : InMux
    port map (
            O => \N__20116\,
            I => \N__20086\
        );

    \I__4557\ : Span4Mux_h
    port map (
            O => \N__20113\,
            I => \N__20083\
        );

    \I__4556\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20078\
        );

    \I__4555\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20078\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20075\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__20101\,
            I => \N__20072\
        );

    \I__4552\ : Span4Mux_v
    port map (
            O => \N__20098\,
            I => \N__20067\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__20089\,
            I => \N__20062\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__20086\,
            I => \N__20062\
        );

    \I__4549\ : Span4Mux_h
    port map (
            O => \N__20083\,
            I => \N__20059\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20052\
        );

    \I__4547\ : Span4Mux_h
    port map (
            O => \N__20075\,
            I => \N__20052\
        );

    \I__4546\ : Span4Mux_h
    port map (
            O => \N__20072\,
            I => \N__20052\
        );

    \I__4545\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20049\
        );

    \I__4544\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20046\
        );

    \I__4543\ : Odrv4
    port map (
            O => \N__20067\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__4542\ : Odrv4
    port map (
            O => \N__20062\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__20059\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__20052\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__20049\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__20046\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\
        );

    \I__4537\ : InMux
    port map (
            O => \N__20033\,
            I => \N__20028\
        );

    \I__4536\ : InMux
    port map (
            O => \N__20032\,
            I => \N__20021\
        );

    \I__4535\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20021\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__20028\,
            I => \N__20015\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__20027\,
            I => \N__20011\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__20026\,
            I => \N__20008\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__20021\,
            I => \N__20005\
        );

    \I__4530\ : InMux
    port map (
            O => \N__20020\,
            I => \N__20002\
        );

    \I__4529\ : InMux
    port map (
            O => \N__20019\,
            I => \N__19997\
        );

    \I__4528\ : InMux
    port map (
            O => \N__20018\,
            I => \N__19997\
        );

    \I__4527\ : Span4Mux_v
    port map (
            O => \N__20015\,
            I => \N__19993\
        );

    \I__4526\ : InMux
    port map (
            O => \N__20014\,
            I => \N__19986\
        );

    \I__4525\ : InMux
    port map (
            O => \N__20011\,
            I => \N__19986\
        );

    \I__4524\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19986\
        );

    \I__4523\ : Span4Mux_h
    port map (
            O => \N__20005\,
            I => \N__19983\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19978\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__19997\,
            I => \N__19978\
        );

    \I__4520\ : InMux
    port map (
            O => \N__19996\,
            I => \N__19975\
        );

    \I__4519\ : Sp12to4
    port map (
            O => \N__19993\,
            I => \N__19970\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__19986\,
            I => \N__19970\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__19983\,
            I => measured_delay_tr_15
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__19978\,
            I => measured_delay_tr_15
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__19975\,
            I => measured_delay_tr_15
        );

    \I__4514\ : Odrv12
    port map (
            O => \N__19970\,
            I => measured_delay_tr_15
        );

    \I__4513\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__19952\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__4509\ : CEMux
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19946\,
            I => \N__19941\
        );

    \I__4507\ : CEMux
    port map (
            O => \N__19945\,
            I => \N__19938\
        );

    \I__4506\ : CEMux
    port map (
            O => \N__19944\,
            I => \N__19935\
        );

    \I__4505\ : Span4Mux_v
    port map (
            O => \N__19941\,
            I => \N__19930\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__19938\,
            I => \N__19930\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19926\
        );

    \I__4502\ : Span4Mux_h
    port map (
            O => \N__19930\,
            I => \N__19923\
        );

    \I__4501\ : CEMux
    port map (
            O => \N__19929\,
            I => \N__19920\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__19926\,
            I => \N__19917\
        );

    \I__4499\ : Span4Mux_h
    port map (
            O => \N__19923\,
            I => \N__19914\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__19920\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__4497\ : Odrv4
    port map (
            O => \N__19917\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__19914\,
            I => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__4495\ : CascadeMux
    port map (
            O => \N__19907\,
            I => \N__19895\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19888\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__19905\,
            I => \N__19885\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19882\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__19903\,
            I => \N__19879\
        );

    \I__4490\ : CascadeMux
    port map (
            O => \N__19902\,
            I => \N__19874\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__19901\,
            I => \N__19870\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__19900\,
            I => \N__19867\
        );

    \I__4487\ : CascadeMux
    port map (
            O => \N__19899\,
            I => \N__19864\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__19898\,
            I => \N__19861\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19854\
        );

    \I__4484\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19837\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19837\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19837\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19837\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19837\
        );

    \I__4479\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19837\
        );

    \I__4478\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19837\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19837\
        );

    \I__4476\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19830\
        );

    \I__4475\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19830\
        );

    \I__4474\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19830\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__19873\,
            I => \N__19827\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19810\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19810\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19810\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19861\,
            I => \N__19810\
        );

    \I__4468\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19810\
        );

    \I__4467\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19810\
        );

    \I__4466\ : InMux
    port map (
            O => \N__19858\,
            I => \N__19810\
        );

    \I__4465\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19810\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19807\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__19837\,
            I => \N__19802\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__19830\,
            I => \N__19802\
        );

    \I__4461\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19799\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19794\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__19807\,
            I => \N__19794\
        );

    \I__4458\ : Span4Mux_v
    port map (
            O => \N__19802\,
            I => \N__19791\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19785\
        );

    \I__4456\ : Sp12to4
    port map (
            O => \N__19794\,
            I => \N__19782\
        );

    \I__4455\ : Span4Mux_h
    port map (
            O => \N__19791\,
            I => \N__19779\
        );

    \I__4454\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19776\
        );

    \I__4453\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19773\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19770\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__19785\,
            I => \N__19767\
        );

    \I__4450\ : Span12Mux_s5_h
    port map (
            O => \N__19782\,
            I => \N__19758\
        );

    \I__4449\ : Sp12to4
    port map (
            O => \N__19779\,
            I => \N__19758\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19776\,
            I => \N__19758\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__19773\,
            I => \N__19758\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__19770\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__4445\ : Odrv4
    port map (
            O => \N__19767\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__4444\ : Odrv12
    port map (
            O => \N__19758\,
            I => \phase_controller_slave.start_timer_trZ0\
        );

    \I__4443\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__4441\ : Odrv4
    port map (
            O => \N__19745\,
            I => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__19736\,
            I => \N__19731\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19728\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19725\
        );

    \I__4435\ : Odrv12
    port map (
            O => \N__19731\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__19728\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__19725\,
            I => \phase_controller_inst1.stoper_tr.time_passed11\
        );

    \I__4432\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19710\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19707\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19702\
        );

    \I__4428\ : Span4Mux_h
    port map (
            O => \N__19710\,
            I => \N__19697\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19707\,
            I => \N__19697\
        );

    \I__4426\ : InMux
    port map (
            O => \N__19706\,
            I => \N__19692\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19705\,
            I => \N__19692\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19702\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__4423\ : Odrv4
    port map (
            O => \N__19697\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__19692\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__4421\ : CascadeMux
    port map (
            O => \N__19685\,
            I => \N__19680\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \N__19677\
        );

    \I__4419\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19674\
        );

    \I__4418\ : InMux
    port map (
            O => \N__19680\,
            I => \N__19669\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19669\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__19674\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19669\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19664\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__19661\,
            I => \N__19656\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__19660\,
            I => \N__19653\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19650\
        );

    \I__4410\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19645\
        );

    \I__4409\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19645\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19650\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19645\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19640\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__4405\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19632\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19629\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19635\,
            I => \N__19626\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19623\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__19629\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19626\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__19623\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19616\,
            I => \bfn_9_29_0_\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19608\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19605\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19602\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19608\,
            I => \N__19599\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__19605\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19602\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__19599\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19592\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__19589\,
            I => \N__19584\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__19588\,
            I => \N__19581\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19578\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19584\,
            I => \N__19573\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19581\,
            I => \N__19573\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19578\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19573\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19568\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__19565\,
            I => \N__19560\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__19564\,
            I => \N__19557\
        );

    \I__4379\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19554\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19549\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19549\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19554\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__19549\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19544\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19537\
        );

    \I__4372\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19534\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19537\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__19534\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19529\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19526\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19519\
        );

    \I__4366\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19516\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19519\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19516\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__4363\ : IoInMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__4361\ : Span12Mux_s6_v
    port map (
            O => \N__19505\,
            I => \N__19502\
        );

    \I__4360\ : Span12Mux_v
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__4359\ : Odrv12
    port map (
            O => \N__19499\,
            I => \delay_measurement_inst.delay_tr_timer.N_138_i\
        );

    \I__4358\ : CascadeMux
    port map (
            O => \N__19496\,
            I => \N__19491\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__19495\,
            I => \N__19488\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19485\
        );

    \I__4355\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19480\
        );

    \I__4354\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19480\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__19485\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__19480\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19475\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__19472\,
            I => \N__19467\
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__19471\,
            I => \N__19464\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19461\
        );

    \I__4347\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19456\
        );

    \I__4346\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19456\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__19461\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__19456\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19451\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19443\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19440\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19437\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19443\,
            I => \N__19434\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__19440\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__19437\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__19434\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__4335\ : InMux
    port map (
            O => \N__19427\,
            I => \bfn_9_28_0_\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19419\
        );

    \I__4333\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19416\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19413\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19419\,
            I => \N__19410\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19416\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19413\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__19410\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19403\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__4326\ : CascadeMux
    port map (
            O => \N__19400\,
            I => \N__19395\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__19399\,
            I => \N__19392\
        );

    \I__4324\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19389\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19395\,
            I => \N__19384\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19392\,
            I => \N__19384\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19389\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19384\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__4319\ : InMux
    port map (
            O => \N__19379\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__19376\,
            I => \N__19371\
        );

    \I__4317\ : CascadeMux
    port map (
            O => \N__19375\,
            I => \N__19368\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19365\
        );

    \I__4315\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19360\
        );

    \I__4314\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19360\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19365\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__19360\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__4311\ : InMux
    port map (
            O => \N__19355\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19347\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19342\
        );

    \I__4308\ : InMux
    port map (
            O => \N__19350\,
            I => \N__19342\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__19347\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__19342\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19337\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19329\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19324\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19324\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19329\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19324\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__4299\ : InMux
    port map (
            O => \N__19319\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19311\
        );

    \I__4297\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19306\
        );

    \I__4296\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19306\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__19311\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__19306\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__4293\ : InMux
    port map (
            O => \N__19301\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__4292\ : CascadeMux
    port map (
            O => \N__19298\,
            I => \N__19293\
        );

    \I__4291\ : CascadeMux
    port map (
            O => \N__19297\,
            I => \N__19290\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19287\
        );

    \I__4289\ : InMux
    port map (
            O => \N__19293\,
            I => \N__19282\
        );

    \I__4288\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19282\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__19287\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19282\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19277\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__19274\,
            I => \N__19269\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__19273\,
            I => \N__19266\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19263\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19258\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19258\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19263\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19258\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__4277\ : InMux
    port map (
            O => \N__19253\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19245\
        );

    \I__4275\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19242\
        );

    \I__4274\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19239\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__19245\,
            I => \N__19236\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19242\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__19239\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__19236\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__4269\ : InMux
    port map (
            O => \N__19229\,
            I => \bfn_9_27_0_\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19221\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19218\
        );

    \I__4266\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19215\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__19221\,
            I => \N__19212\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__19218\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__19215\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__19212\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__4261\ : InMux
    port map (
            O => \N__19205\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__4260\ : CascadeMux
    port map (
            O => \N__19202\,
            I => \N__19197\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__19201\,
            I => \N__19194\
        );

    \I__4258\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19191\
        );

    \I__4257\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19186\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19186\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__19191\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__19186\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19181\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__19178\,
            I => \N__19173\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__19177\,
            I => \N__19170\
        );

    \I__4250\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19167\
        );

    \I__4249\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19162\
        );

    \I__4248\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19162\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__19167\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__19162\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__4245\ : InMux
    port map (
            O => \N__19157\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__4244\ : InMux
    port map (
            O => \N__19154\,
            I => \N__19149\
        );

    \I__4243\ : InMux
    port map (
            O => \N__19153\,
            I => \N__19144\
        );

    \I__4242\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19144\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__19149\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__19144\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__4239\ : InMux
    port map (
            O => \N__19139\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__4238\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19131\
        );

    \I__4237\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19126\
        );

    \I__4236\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19126\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__19131\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__19126\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__4233\ : InMux
    port map (
            O => \N__19121\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__19118\,
            I => \N__19089\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__19117\,
            I => \N__19085\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__19116\,
            I => \N__19082\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__19115\,
            I => \N__19078\
        );

    \I__4228\ : CascadeMux
    port map (
            O => \N__19114\,
            I => \N__19074\
        );

    \I__4227\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19055\
        );

    \I__4226\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19055\
        );

    \I__4225\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19055\
        );

    \I__4224\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19055\
        );

    \I__4223\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19055\
        );

    \I__4222\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19055\
        );

    \I__4221\ : InMux
    port map (
            O => \N__19107\,
            I => \N__19055\
        );

    \I__4220\ : InMux
    port map (
            O => \N__19106\,
            I => \N__19055\
        );

    \I__4219\ : InMux
    port map (
            O => \N__19105\,
            I => \N__19038\
        );

    \I__4218\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19038\
        );

    \I__4217\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19038\
        );

    \I__4216\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19038\
        );

    \I__4215\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19038\
        );

    \I__4214\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19038\
        );

    \I__4213\ : InMux
    port map (
            O => \N__19099\,
            I => \N__19038\
        );

    \I__4212\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19038\
        );

    \I__4211\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19021\
        );

    \I__4210\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19021\
        );

    \I__4209\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19021\
        );

    \I__4208\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19021\
        );

    \I__4207\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19021\
        );

    \I__4206\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19021\
        );

    \I__4205\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19021\
        );

    \I__4204\ : InMux
    port map (
            O => \N__19088\,
            I => \N__19021\
        );

    \I__4203\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19004\
        );

    \I__4202\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19004\
        );

    \I__4201\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19004\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19004\
        );

    \I__4199\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19004\
        );

    \I__4198\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19004\
        );

    \I__4197\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19004\
        );

    \I__4196\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19004\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__19055\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__19038\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__19021\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__19004\,
            I => \delay_measurement_inst.un1_elapsed_time_hc\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18965\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18965\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18965\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18965\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18965\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18965\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18954\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18954\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18954\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18986\,
            I => \N__18954\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18954\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18984\,
            I => \N__18949\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18949\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18938\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18938\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18938\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18938\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18938\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__18965\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__18954\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__18949\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__18938\,
            I => \delay_measurement_inst.delay_hc_reg3lto31_0_0\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \N__18925\
        );

    \I__4168\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18922\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18919\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18922\,
            I => measured_delay_hc_26
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__18919\,
            I => measured_delay_hc_26
        );

    \I__4164\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18911\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__18911\,
            I => \N__18908\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__18908\,
            I => \N__18904\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__4160\ : Odrv4
    port map (
            O => \N__18904\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18901\,
            I => \delay_measurement_inst.elapsed_time_hc_1\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18889\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__18892\,
            I => \N__18885\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18889\,
            I => \N__18882\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18879\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18876\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__18882\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18879\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__18876\,
            I => \delay_measurement_inst.elapsed_time_hc_2\
        );

    \I__4149\ : CEMux
    port map (
            O => \N__18869\,
            I => \N__18854\
        );

    \I__4148\ : CEMux
    port map (
            O => \N__18868\,
            I => \N__18854\
        );

    \I__4147\ : CEMux
    port map (
            O => \N__18867\,
            I => \N__18854\
        );

    \I__4146\ : CEMux
    port map (
            O => \N__18866\,
            I => \N__18854\
        );

    \I__4145\ : CEMux
    port map (
            O => \N__18865\,
            I => \N__18854\
        );

    \I__4144\ : GlobalMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__4143\ : gio2CtrlBuf
    port map (
            O => \N__18851\,
            I => \delay_measurement_inst.delay_hc_timer.N_136_i_g\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18843\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18840\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18837\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18843\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18840\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18837\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18830\,
            I => \bfn_9_26_0_\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18822\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18819\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18825\,
            I => \N__18816\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__18822\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18819\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__18816\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18809\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__18806\,
            I => \N__18801\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18805\,
            I => \N__18798\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18795\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18790\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18790\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18795\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__18790\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18785\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__18782\,
            I => \N__18777\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__18781\,
            I => \N__18774\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18771\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18766\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18766\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18771\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__18766\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__4113\ : InMux
    port map (
            O => \N__18761\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18753\
        );

    \I__4111\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18748\
        );

    \I__4110\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18748\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__18753\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__18748\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18743\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18732\
        );

    \I__4104\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18729\
        );

    \I__4103\ : InMux
    port map (
            O => \N__18735\,
            I => \N__18726\
        );

    \I__4102\ : Span4Mux_v
    port map (
            O => \N__18732\,
            I => \N__18721\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18729\,
            I => \N__18721\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18718\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__18721\,
            I => \N__18715\
        );

    \I__4098\ : Odrv12
    port map (
            O => \N__18718\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__18715\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18706\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__18709\,
            I => \N__18703\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__4093\ : InMux
    port map (
            O => \N__18703\,
            I => \N__18697\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__18700\,
            I => \N__18692\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__18697\,
            I => \N__18692\
        );

    \I__4090\ : Span4Mux_h
    port map (
            O => \N__18692\,
            I => \N__18688\
        );

    \I__4089\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18685\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__18688\,
            I => \N__18682\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18685\,
            I => \N__18679\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__18682\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\
        );

    \I__4085\ : Odrv12
    port map (
            O => \N__18679\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__18674\,
            I => \N__18670\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__4082\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__18667\,
            I => measured_delay_hc_30
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18664\,
            I => measured_delay_hc_30
        );

    \I__4079\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18655\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18652\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__18655\,
            I => measured_delay_hc_24
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__18652\,
            I => measured_delay_hc_24
        );

    \I__4075\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18643\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18640\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__18643\,
            I => measured_delay_hc_25
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__18640\,
            I => measured_delay_hc_25
        );

    \I__4071\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18631\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18628\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__18631\,
            I => measured_delay_hc_28
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18628\,
            I => measured_delay_hc_28
        );

    \I__4067\ : InMux
    port map (
            O => \N__18623\,
            I => \N__18619\
        );

    \I__4066\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18616\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__18619\,
            I => measured_delay_hc_29
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__18616\,
            I => measured_delay_hc_29
        );

    \I__4063\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18593\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18593\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18586\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18608\,
            I => \N__18586\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18586\
        );

    \I__4058\ : InMux
    port map (
            O => \N__18606\,
            I => \N__18573\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18573\
        );

    \I__4056\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18573\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18573\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18573\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18573\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18566\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18566\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18566\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__18593\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__18586\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__18573\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__18566\,
            I => \delay_measurement_inst.delay_hc_reg3\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18553\
        );

    \I__4044\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18550\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__18553\,
            I => measured_delay_hc_23
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18550\,
            I => measured_delay_hc_23
        );

    \I__4041\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18541\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18538\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__18541\,
            I => measured_delay_hc_27
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18538\,
            I => measured_delay_hc_27
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__18527\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18524\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__4033\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18517\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18514\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__18517\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__18514\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18509\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__18503\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\
        );

    \I__4026\ : CEMux
    port map (
            O => \N__18500\,
            I => \N__18496\
        );

    \I__4025\ : CEMux
    port map (
            O => \N__18499\,
            I => \N__18493\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__18496\,
            I => \N__18488\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__18493\,
            I => \N__18484\
        );

    \I__4022\ : CEMux
    port map (
            O => \N__18492\,
            I => \N__18481\
        );

    \I__4021\ : CEMux
    port map (
            O => \N__18491\,
            I => \N__18478\
        );

    \I__4020\ : Span4Mux_v
    port map (
            O => \N__18488\,
            I => \N__18475\
        );

    \I__4019\ : CEMux
    port map (
            O => \N__18487\,
            I => \N__18472\
        );

    \I__4018\ : Span4Mux_h
    port map (
            O => \N__18484\,
            I => \N__18467\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18467\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__18478\,
            I => \N__18464\
        );

    \I__4015\ : Span4Mux_h
    port map (
            O => \N__18475\,
            I => \N__18459\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18472\,
            I => \N__18459\
        );

    \I__4013\ : Sp12to4
    port map (
            O => \N__18467\,
            I => \N__18456\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__18464\,
            I => \N__18451\
        );

    \I__4011\ : Span4Mux_h
    port map (
            O => \N__18459\,
            I => \N__18451\
        );

    \I__4010\ : Odrv12
    port map (
            O => \N__18456\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__18451\,
            I => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18443\,
            I => \N__18439\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18442\,
            I => \N__18435\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__18439\,
            I => \N__18432\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18429\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__18435\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__18432\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__18429\,
            I => \phase_controller_inst1.stoper_hc.time_passed11\
        );

    \I__4000\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18415\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18418\,
            I => \N__18411\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__18415\,
            I => \N__18408\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18405\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18411\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__18408\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18405\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__18395\,
            I => \N__18389\
        );

    \I__3990\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18384\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18393\,
            I => \N__18379\
        );

    \I__3988\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18379\
        );

    \I__3987\ : Span4Mux_h
    port map (
            O => \N__18389\,
            I => \N__18376\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18371\
        );

    \I__3985\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18371\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__18384\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__18379\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__18376\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__18371\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18359\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__3978\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18353\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__18353\,
            I => \phase_controller_slave.start_timer_hc_0_sqmuxa\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__18350\,
            I => \N__18344\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__18349\,
            I => \N__18341\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__18348\,
            I => \N__18338\
        );

    \I__3973\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18318\
        );

    \I__3972\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18309\
        );

    \I__3971\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18309\
        );

    \I__3970\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18309\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18302\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18336\,
            I => \N__18302\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18302\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18285\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18285\
        );

    \I__3964\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18285\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18285\
        );

    \I__3962\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18285\
        );

    \I__3961\ : InMux
    port map (
            O => \N__18329\,
            I => \N__18285\
        );

    \I__3960\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18285\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18285\
        );

    \I__3958\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18274\
        );

    \I__3957\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18274\
        );

    \I__3956\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18274\
        );

    \I__3955\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18274\
        );

    \I__3954\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18274\
        );

    \I__3953\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18271\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__18318\,
            I => \N__18268\
        );

    \I__3951\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18262\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18262\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__18309\,
            I => \N__18255\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__18302\,
            I => \N__18255\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18255\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N__18248\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18248\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__18268\,
            I => \N__18248\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18267\,
            I => \N__18245\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__18262\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3941\ : Odrv12
    port map (
            O => \N__18255\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__18248\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__18245\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18212\
        );

    \I__3937\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18198\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18198\
        );

    \I__3935\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18198\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18198\
        );

    \I__3933\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18198\
        );

    \I__3932\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18198\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18181\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18181\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18181\
        );

    \I__3928\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18181\
        );

    \I__3927\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18181\
        );

    \I__3926\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18181\
        );

    \I__3925\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18181\
        );

    \I__3924\ : InMux
    port map (
            O => \N__18222\,
            I => \N__18181\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18170\
        );

    \I__3922\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18170\
        );

    \I__3921\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18170\
        );

    \I__3920\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18170\
        );

    \I__3919\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18170\
        );

    \I__3918\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18167\
        );

    \I__3917\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18164\
        );

    \I__3916\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18158\
        );

    \I__3915\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18158\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__18198\,
            I => \N__18155\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__18181\,
            I => \N__18146\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__18170\,
            I => \N__18146\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__18167\,
            I => \N__18146\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__18164\,
            I => \N__18146\
        );

    \I__3909\ : InMux
    port map (
            O => \N__18163\,
            I => \N__18143\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__18158\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3907\ : Odrv12
    port map (
            O => \N__18155\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__18146\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__18143\,
            I => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__3903\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__18128\,
            I => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__3901\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__18122\,
            I => \phase_controller_slave.N_21\
        );

    \I__3899\ : IoInMux
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18116\,
            I => \N__18113\
        );

    \I__3897\ : Odrv12
    port map (
            O => \N__18113\,
            I => s3_phy_c
        );

    \I__3896\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18106\
        );

    \I__3895\ : CascadeMux
    port map (
            O => \N__18109\,
            I => \N__18103\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__18106\,
            I => \N__18098\
        );

    \I__3893\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18091\
        );

    \I__3892\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18091\
        );

    \I__3891\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18091\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__18098\,
            I => \N__18088\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__18091\,
            I => \N__18085\
        );

    \I__3888\ : Span4Mux_h
    port map (
            O => \N__18088\,
            I => \N__18080\
        );

    \I__3887\ : Span4Mux_h
    port map (
            O => \N__18085\,
            I => \N__18080\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__18080\,
            I => \phase_controller_slave.stoper_hc.time_passed11\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__3884\ : InMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__18065\,
            I => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\
        );

    \I__3880\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18057\
        );

    \I__3879\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18052\
        );

    \I__3878\ : InMux
    port map (
            O => \N__18060\,
            I => \N__18052\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__18057\,
            I => \N__18047\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__18052\,
            I => \N__18044\
        );

    \I__3875\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18039\
        );

    \I__3874\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18039\
        );

    \I__3873\ : Odrv12
    port map (
            O => \N__18047\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__18044\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__18039\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__3870\ : InMux
    port map (
            O => \N__18032\,
            I => \N__18028\
        );

    \I__3869\ : InMux
    port map (
            O => \N__18031\,
            I => \N__18025\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__18028\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__18025\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__3866\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__18017\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\
        );

    \I__3864\ : InMux
    port map (
            O => \N__18014\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__3863\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18007\
        );

    \I__3862\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18004\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__18007\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__18004\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__17996\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\
        );

    \I__3857\ : InMux
    port map (
            O => \N__17993\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17986\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17983\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17986\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17983\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17975\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17972\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__3849\ : InMux
    port map (
            O => \N__17969\,
            I => \N__17965\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17962\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__17965\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17962\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17954\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__17954\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\
        );

    \I__3843\ : InMux
    port map (
            O => \N__17951\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__3842\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17944\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17941\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17944\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__17941\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__3838\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__17933\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17930\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__3835\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17923\
        );

    \I__3834\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17920\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__17923\,
            I => \N__17917\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17920\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__17917\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17909\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\
        );

    \I__3828\ : InMux
    port map (
            O => \N__17906\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17899\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17896\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__17899\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__17896\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__17891\,
            I => \N__17888\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17885\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__17885\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\
        );

    \I__3820\ : InMux
    port map (
            O => \N__17882\,
            I => \bfn_9_19_0_\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17875\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17878\,
            I => \N__17872\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__17875\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__17872\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17863\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17860\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17863\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17860\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__3810\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17849\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__17840\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\
        );

    \I__3805\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__17834\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17831\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17824\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17821\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__17824\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__17821\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17813\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17810\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17803\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17800\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__17803\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__17800\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__17792\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17789\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17782\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17779\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17782\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17779\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17771\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\
        );

    \I__3782\ : InMux
    port map (
            O => \N__17768\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17761\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17764\,
            I => \N__17758\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__17761\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17758\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__17750\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17747\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17741\,
            I => \N__17738\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__17738\,
            I => \N__17734\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17731\
        );

    \I__3770\ : Odrv4
    port map (
            O => \N__17734\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__17731\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__17726\,
            I => \N__17723\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__17717\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\
        );

    \I__3764\ : InMux
    port map (
            O => \N__17714\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__3763\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17707\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17704\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__17707\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__17704\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__17696\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17693\,
            I => \bfn_9_18_0_\
        );

    \I__3756\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17686\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17689\,
            I => \N__17683\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__17686\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__17683\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__3752\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__17675\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\
        );

    \I__3750\ : InMux
    port map (
            O => \N__17672\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__3749\ : InMux
    port map (
            O => \N__17669\,
            I => \N__17665\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17662\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__17665\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__17662\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17651\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17651\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17648\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__3741\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17641\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17638\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17641\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17638\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__17630\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17627\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17620\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17617\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__17620\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17617\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17609\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\
        );

    \I__3728\ : InMux
    port map (
            O => \N__17606\,
            I => \bfn_9_15_0_\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17599\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17596\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17599\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__17596\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__17588\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17585\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17578\
        );

    \I__3719\ : InMux
    port map (
            O => \N__17581\,
            I => \N__17575\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17578\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__17575\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17570\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__17564\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \N__17553\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__17560\,
            I => \N__17550\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__17559\,
            I => \N__17547\
        );

    \I__3710\ : CascadeMux
    port map (
            O => \N__17558\,
            I => \N__17544\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__17557\,
            I => \N__17536\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__17556\,
            I => \N__17533\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17516\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17516\
        );

    \I__3705\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17516\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17516\
        );

    \I__3703\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17509\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17509\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17509\
        );

    \I__3700\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17501\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17501\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17496\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17496\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17479\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17479\
        );

    \I__3694\ : InMux
    port map (
            O => \N__17530\,
            I => \N__17479\
        );

    \I__3693\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17479\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17528\,
            I => \N__17479\
        );

    \I__3691\ : InMux
    port map (
            O => \N__17527\,
            I => \N__17479\
        );

    \I__3690\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17479\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17479\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__17516\,
            I => \N__17474\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17509\,
            I => \N__17474\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__17508\,
            I => \N__17471\
        );

    \I__3685\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17466\
        );

    \I__3684\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17463\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17501\,
            I => \N__17460\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__17496\,
            I => \N__17453\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__17479\,
            I => \N__17453\
        );

    \I__3680\ : Span4Mux_h
    port map (
            O => \N__17474\,
            I => \N__17453\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17446\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17470\,
            I => \N__17446\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17469\,
            I => \N__17446\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17466\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__17463\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__17460\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3673\ : Odrv4
    port map (
            O => \N__17453\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__17446\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__3671\ : CascadeMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17422\
        );

    \I__3669\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17407\
        );

    \I__3668\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17407\
        );

    \I__3667\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17407\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17407\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17427\,
            I => \N__17407\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17407\
        );

    \I__3663\ : InMux
    port map (
            O => \N__17425\,
            I => \N__17407\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__17422\,
            I => \N__17391\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__17407\,
            I => \N__17388\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17406\,
            I => \N__17373\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17405\,
            I => \N__17373\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17373\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17403\,
            I => \N__17373\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17402\,
            I => \N__17373\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17373\
        );

    \I__3654\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17373\
        );

    \I__3653\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17367\
        );

    \I__3652\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17364\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17355\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17355\
        );

    \I__3649\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17355\
        );

    \I__3648\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17355\
        );

    \I__3647\ : Span4Mux_v
    port map (
            O => \N__17391\,
            I => \N__17352\
        );

    \I__3646\ : Span4Mux_h
    port map (
            O => \N__17388\,
            I => \N__17347\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__17373\,
            I => \N__17347\
        );

    \I__3644\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17340\
        );

    \I__3643\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17340\
        );

    \I__3642\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17340\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__17367\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__17364\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17355\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3638\ : Odrv4
    port map (
            O => \N__17352\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__17347\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__17340\,
            I => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__3634\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__17321\,
            I => \N__17318\
        );

    \I__3632\ : Span4Mux_h
    port map (
            O => \N__17318\,
            I => \N__17315\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__17315\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17312\,
            I => \N__17308\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17305\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17308\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__17305\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17297\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17297\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17294\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__3623\ : InMux
    port map (
            O => \N__17291\,
            I => \N__17287\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17290\,
            I => \N__17284\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__17287\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__17284\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__3619\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__17276\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\
        );

    \I__3617\ : InMux
    port map (
            O => \N__17273\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__3616\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17266\
        );

    \I__3615\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17263\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__17266\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__17263\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__3612\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17255\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\
        );

    \I__3610\ : InMux
    port map (
            O => \N__17252\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__3609\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17245\
        );

    \I__3608\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17242\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__17245\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__17242\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__3605\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17234\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__17234\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\
        );

    \I__3603\ : InMux
    port map (
            O => \N__17231\,
            I => \bfn_9_14_0_\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17228\,
            I => \N__17224\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17221\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__17224\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__17221\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17213\,
            I => \N__17210\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__17210\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\
        );

    \I__3595\ : InMux
    port map (
            O => \N__17207\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__3594\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17200\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17197\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__17200\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__17197\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__3590\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__17189\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\
        );

    \I__3588\ : InMux
    port map (
            O => \N__17186\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__3587\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__17180\,
            I => \N__17176\
        );

    \I__3585\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__3584\ : Span4Mux_h
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__17173\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__17170\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__3581\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17162\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__17162\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\
        );

    \I__3579\ : InMux
    port map (
            O => \N__17159\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__3578\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17152\
        );

    \I__3577\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__17152\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__17149\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__3573\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17138\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__17138\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\
        );

    \I__3571\ : InMux
    port map (
            O => \N__17135\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__3570\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17128\
        );

    \I__3569\ : InMux
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__17128\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__17125\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__3566\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__17117\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\
        );

    \I__3564\ : InMux
    port map (
            O => \N__17114\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__3562\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__17105\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__3560\ : InMux
    port map (
            O => \N__17102\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__3559\ : InMux
    port map (
            O => \N__17099\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__17096\,
            I => \N__17092\
        );

    \I__3557\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17087\
        );

    \I__3556\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17087\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__17087\,
            I => \N__17084\
        );

    \I__3554\ : Span4Mux_v
    port map (
            O => \N__17084\,
            I => \N__17080\
        );

    \I__3553\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__17080\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__17077\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__3550\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17068\
        );

    \I__3549\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17064\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17061\
        );

    \I__3547\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17058\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__17064\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__17061\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__17058\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__3542\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__17039\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\
        );

    \I__3538\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17032\
        );

    \I__3537\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__17032\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__17029\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__3534\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__17021\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\
        );

    \I__3532\ : InMux
    port map (
            O => \N__17018\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__3531\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17011\
        );

    \I__3530\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17008\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__17011\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__17008\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__3526\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__16994\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16988\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16985\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16978\
        );

    \I__3519\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16975\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__16978\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__16975\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16967\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\
        );

    \I__3514\ : InMux
    port map (
            O => \N__16964\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16957\
        );

    \I__3512\ : InMux
    port map (
            O => \N__16960\,
            I => \N__16954\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__16957\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__16954\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__3509\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16946\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16946\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16943\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16940\,
            I => \N__16936\
        );

    \I__3505\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16933\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16936\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__16933\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16925\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16925\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16922\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \N__16916\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16910\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16910\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__16910\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__3495\ : InMux
    port map (
            O => \N__16907\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__16901\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16898\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__16892\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16889\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__16883\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16880\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \N__16874\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16871\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16871\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__3482\ : InMux
    port map (
            O => \N__16868\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__3481\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16862\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16862\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16859\,
            I => \bfn_8_29_0_\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16853\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__16853\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16850\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__3475\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__16844\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16841\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16835\,
            I => \N__16829\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16826\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16823\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16820\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16829\,
            I => \N__16813\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16826\,
            I => \N__16813\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__16823\,
            I => \N__16813\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__16820\,
            I => \N__16810\
        );

    \I__3463\ : Span4Mux_v
    port map (
            O => \N__16813\,
            I => \N__16807\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__16810\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__16807\,
            I => \delay_measurement_inst.delay_hc_reg3lto14\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16802\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__16799\,
            I => \N__16789\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16798\,
            I => \N__16786\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16797\,
            I => \N__16783\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16774\
        );

    \I__3455\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16774\
        );

    \I__3454\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16774\
        );

    \I__3453\ : InMux
    port map (
            O => \N__16793\,
            I => \N__16774\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16792\,
            I => \N__16769\
        );

    \I__3451\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16769\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__16786\,
            I => \N__16762\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__16783\,
            I => \N__16762\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__16774\,
            I => \N__16762\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__16769\,
            I => \N__16759\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__16762\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__16759\,
            I => \delay_measurement_inst.delay_hc_reg3lto15\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16754\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__16751\,
            I => \N__16748\
        );

    \I__3442\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16743\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16740\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__16746\,
            I => \N__16737\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__16743\,
            I => \N__16732\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__16740\,
            I => \N__16732\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16729\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__16732\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__16729\,
            I => \delay_measurement_inst.elapsed_time_hc_16\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16724\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16714\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16711\
        );

    \I__3430\ : Span4Mux_h
    port map (
            O => \N__16714\,
            I => \N__16705\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__16711\,
            I => \N__16705\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16702\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__16705\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__16702\,
            I => \delay_measurement_inst.elapsed_time_hc_17\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16697\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__16691\,
            I => \N__16687\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16684\
        );

    \I__3421\ : Span4Mux_h
    port map (
            O => \N__16687\,
            I => \N__16678\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16684\,
            I => \N__16678\
        );

    \I__3419\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16675\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__16678\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16675\,
            I => \delay_measurement_inst.elapsed_time_hc_18\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16670\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16663\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__16666\,
            I => \N__16659\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__16663\,
            I => \N__16656\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16653\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16650\
        );

    \I__3410\ : Span4Mux_h
    port map (
            O => \N__16656\,
            I => \N__16643\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__16653\,
            I => \N__16643\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16650\,
            I => \N__16643\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__16643\,
            I => \delay_measurement_inst.elapsed_time_hc_19\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16640\,
            I => \bfn_8_28_0_\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16630\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16627\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__16630\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16627\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16622\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16613\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16613\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__16613\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16610\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__16607\,
            I => \N__16603\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16606\,
            I => \N__16600\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16597\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16600\,
            I => \N__16593\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__16597\,
            I => \N__16590\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16587\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__16593\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__16590\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__16587\,
            I => \delay_measurement_inst.elapsed_time_hc_5\
        );

    \I__3386\ : InMux
    port map (
            O => \N__16580\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3385\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16574\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__16574\,
            I => \N__16569\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16566\
        );

    \I__3382\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16563\
        );

    \I__3381\ : Odrv4
    port map (
            O => \N__16569\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__16566\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16563\,
            I => \delay_measurement_inst.delay_hc_reg3lto6\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16556\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3377\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16550\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16550\,
            I => \N__16545\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16540\
        );

    \I__3374\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16540\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__16545\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16540\,
            I => \delay_measurement_inst.elapsed_time_hc_7\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16535\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16532\,
            I => \N__16528\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__16531\,
            I => \N__16525\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__16528\,
            I => \N__16521\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16525\,
            I => \N__16516\
        );

    \I__3366\ : InMux
    port map (
            O => \N__16524\,
            I => \N__16516\
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__16521\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__16516\,
            I => \delay_measurement_inst.elapsed_time_hc_8\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16511\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__16508\,
            I => \N__16504\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16500\
        );

    \I__3360\ : InMux
    port map (
            O => \N__16504\,
            I => \N__16497\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16503\,
            I => \N__16494\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16500\,
            I => \N__16490\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__16497\,
            I => \N__16485\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16485\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16482\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__16490\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__3353\ : Odrv12
    port map (
            O => \N__16485\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16482\,
            I => \delay_measurement_inst.delay_hc_reg3lto9\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16475\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3350\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16469\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__16469\,
            I => \N__16464\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16459\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16459\
        );

    \I__3346\ : Odrv12
    port map (
            O => \N__16464\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16459\,
            I => \delay_measurement_inst.elapsed_time_hc_10\
        );

    \I__3344\ : InMux
    port map (
            O => \N__16454\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16446\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16441\
        );

    \I__3341\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16441\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16438\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__16441\,
            I => \N__16435\
        );

    \I__3338\ : Odrv12
    port map (
            O => \N__16438\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__16435\,
            I => \delay_measurement_inst.elapsed_time_hc_11\
        );

    \I__3336\ : InMux
    port map (
            O => \N__16430\,
            I => \bfn_8_27_0_\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16427\,
            I => \N__16422\
        );

    \I__3334\ : InMux
    port map (
            O => \N__16426\,
            I => \N__16419\
        );

    \I__3333\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16416\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16422\,
            I => \N__16413\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__16419\,
            I => \N__16408\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16416\,
            I => \N__16408\
        );

    \I__3329\ : Odrv12
    port map (
            O => \N__16413\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3328\ : Odrv12
    port map (
            O => \N__16408\,
            I => \delay_measurement_inst.elapsed_time_hc_12\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16403\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16396\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__16399\,
            I => \N__16393\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__16396\,
            I => \N__16389\
        );

    \I__3323\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16386\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16392\,
            I => \N__16383\
        );

    \I__3321\ : Span4Mux_h
    port map (
            O => \N__16389\,
            I => \N__16378\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__16386\,
            I => \N__16378\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__16383\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__16378\,
            I => \delay_measurement_inst.elapsed_time_hc_13\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16373\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6_cascade_\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16361\
        );

    \I__3314\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16361\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__16361\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_3\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16358\,
            I => \N__16354\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16351\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__16354\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__16351\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\
        );

    \I__3308\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16339\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16339\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16336\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16339\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16336\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__16328\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__16325\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16322\,
            I => \N__16319\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__16319\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16312\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16315\,
            I => \N__16309\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__16312\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16309\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__16304\,
            I => \N__16301\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16297\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16300\,
            I => \N__16294\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16297\,
            I => \N__16290\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__16294\,
            I => \N__16287\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16284\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__16290\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__16287\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__16284\,
            I => \delay_measurement_inst.elapsed_time_hc_3\
        );

    \I__3285\ : CascadeMux
    port map (
            O => \N__16277\,
            I => \N__16274\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16271\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16271\,
            I => \N__16267\
        );

    \I__3282\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16264\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__16267\,
            I => \N__16258\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__16264\,
            I => \N__16258\
        );

    \I__3279\ : InMux
    port map (
            O => \N__16263\,
            I => \N__16255\
        );

    \I__3278\ : Odrv4
    port map (
            O => \N__16258\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16255\,
            I => \delay_measurement_inst.elapsed_time_hc_4\
        );

    \I__3276\ : InMux
    port map (
            O => \N__16250\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3275\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16244\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1Z0Z_9\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__16241\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_cascade_\
        );

    \I__3272\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16235\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__16235\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__16232\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__16229\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_cascade_\
        );

    \I__3268\ : InMux
    port map (
            O => \N__16226\,
            I => \N__16223\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__16223\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__16220\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_cascade_\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16211\
        );

    \I__3264\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16211\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__16211\,
            I => \N__16208\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__16205\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2\
        );

    \I__3260\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16199\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__16199\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__16196\,
            I => \N__16191\
        );

    \I__3257\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16187\
        );

    \I__3256\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16178\
        );

    \I__3255\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16178\
        );

    \I__3254\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16178\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__16187\,
            I => \N__16175\
        );

    \I__3252\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16172\
        );

    \I__3251\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16169\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__16178\,
            I => \N__16166\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__16175\,
            I => \N__16163\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__16172\,
            I => \N__16160\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__16169\,
            I => \N__16155\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__16166\,
            I => \N__16155\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__16163\,
            I => measured_delay_hc_9
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__16160\,
            I => measured_delay_hc_9
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__16155\,
            I => measured_delay_hc_9
        );

    \I__3242\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16143\
        );

    \I__3241\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16140\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__16146\,
            I => \N__16135\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__16143\,
            I => \N__16130\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__16140\,
            I => \N__16130\
        );

    \I__3237\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16127\
        );

    \I__3236\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16124\
        );

    \I__3235\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16121\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__16130\,
            I => \N__16118\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__16127\,
            I => \N__16113\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__16124\,
            I => \N__16113\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__16121\,
            I => measured_delay_hc_7
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__16118\,
            I => measured_delay_hc_7
        );

    \I__3229\ : Odrv12
    port map (
            O => \N__16113\,
            I => measured_delay_hc_7
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__16106\,
            I => \N__16103\
        );

    \I__3227\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16099\
        );

    \I__3226\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16096\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__16099\,
            I => \N__16090\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__16096\,
            I => \N__16087\
        );

    \I__3223\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16082\
        );

    \I__3222\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16082\
        );

    \I__3221\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16079\
        );

    \I__3220\ : Span4Mux_h
    port map (
            O => \N__16090\,
            I => \N__16076\
        );

    \I__3219\ : Span4Mux_v
    port map (
            O => \N__16087\,
            I => \N__16073\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__16082\,
            I => \N__16070\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__16079\,
            I => measured_delay_hc_2
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__16076\,
            I => measured_delay_hc_2
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__16073\,
            I => measured_delay_hc_2
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__16070\,
            I => measured_delay_hc_2
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__16061\,
            I => \N__16056\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__16060\,
            I => \N__16052\
        );

    \I__3211\ : InMux
    port map (
            O => \N__16059\,
            I => \N__16049\
        );

    \I__3210\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16046\
        );

    \I__3209\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16042\
        );

    \I__3208\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16039\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__16049\,
            I => \N__16036\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__16046\,
            I => \N__16033\
        );

    \I__3205\ : InMux
    port map (
            O => \N__16045\,
            I => \N__16030\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__16042\,
            I => \N__16027\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__16039\,
            I => \N__16018\
        );

    \I__3202\ : Span4Mux_v
    port map (
            O => \N__16036\,
            I => \N__16018\
        );

    \I__3201\ : Span4Mux_h
    port map (
            O => \N__16033\,
            I => \N__16018\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16018\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__16027\,
            I => measured_delay_hc_8
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__16018\,
            I => measured_delay_hc_8
        );

    \I__3197\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__16010\,
            I => \N__16003\
        );

    \I__3195\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16000\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__16008\,
            I => \N__15997\
        );

    \I__3193\ : InMux
    port map (
            O => \N__16007\,
            I => \N__15994\
        );

    \I__3192\ : InMux
    port map (
            O => \N__16006\,
            I => \N__15991\
        );

    \I__3191\ : Span4Mux_v
    port map (
            O => \N__16003\,
            I => \N__15986\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__16000\,
            I => \N__15986\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15983\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__15994\,
            I => \N__15980\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__15991\,
            I => \N__15977\
        );

    \I__3186\ : Span4Mux_h
    port map (
            O => \N__15986\,
            I => \N__15974\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__15983\,
            I => measured_delay_hc_12
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__15980\,
            I => measured_delay_hc_12
        );

    \I__3183\ : Odrv12
    port map (
            O => \N__15977\,
            I => measured_delay_hc_12
        );

    \I__3182\ : Odrv4
    port map (
            O => \N__15974\,
            I => measured_delay_hc_12
        );

    \I__3181\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15962\,
            I => \N__15956\
        );

    \I__3179\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15953\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15949\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15946\
        );

    \I__3176\ : Span4Mux_v
    port map (
            O => \N__15956\,
            I => \N__15941\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__15953\,
            I => \N__15941\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15952\,
            I => \N__15938\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15935\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__15946\,
            I => \N__15932\
        );

    \I__3171\ : Span4Mux_h
    port map (
            O => \N__15941\,
            I => \N__15929\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15938\,
            I => measured_delay_hc_10
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__15935\,
            I => measured_delay_hc_10
        );

    \I__3168\ : Odrv12
    port map (
            O => \N__15932\,
            I => measured_delay_hc_10
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__15929\,
            I => measured_delay_hc_10
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15908\
        );

    \I__3164\ : InMux
    port map (
            O => \N__15916\,
            I => \N__15908\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15908\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__15908\,
            I => \N__15900\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15897\
        );

    \I__3160\ : CascadeMux
    port map (
            O => \N__15906\,
            I => \N__15889\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__15905\,
            I => \N__15886\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15877\
        );

    \I__3157\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15877\
        );

    \I__3156\ : Span4Mux_h
    port map (
            O => \N__15900\,
            I => \N__15866\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__15897\,
            I => \N__15866\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15861\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15861\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15856\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15856\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15847\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15847\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15847\
        );

    \I__3147\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15847\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15884\,
            I => \N__15844\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15839\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15839\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__15877\,
            I => \N__15835\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15824\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15824\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15824\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15873\,
            I => \N__15824\
        );

    \I__3138\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15824\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15821\
        );

    \I__3136\ : Span4Mux_h
    port map (
            O => \N__15866\,
            I => \N__15814\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__15861\,
            I => \N__15814\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15856\,
            I => \N__15814\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15847\,
            I => \N__15807\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15844\,
            I => \N__15807\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__15839\,
            I => \N__15807\
        );

    \I__3130\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15804\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__15835\,
            I => \N__15797\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__15824\,
            I => \N__15797\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__15821\,
            I => \N__15797\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__15814\,
            I => \N__15792\
        );

    \I__3125\ : Span4Mux_v
    port map (
            O => \N__15807\,
            I => \N__15792\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15804\,
            I => measured_delay_hc_31
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__15797\,
            I => measured_delay_hc_31
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__15792\,
            I => measured_delay_hc_31
        );

    \I__3121\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15780\
        );

    \I__3120\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15775\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__15783\,
            I => \N__15772\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__15780\,
            I => \N__15769\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15766\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15763\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__15775\,
            I => \N__15760\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15757\
        );

    \I__3113\ : Span4Mux_h
    port map (
            O => \N__15769\,
            I => \N__15752\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15766\,
            I => \N__15752\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__15763\,
            I => \N__15749\
        );

    \I__3110\ : Span4Mux_h
    port map (
            O => \N__15760\,
            I => \N__15746\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15757\,
            I => measured_delay_hc_11
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__15752\,
            I => measured_delay_hc_11
        );

    \I__3107\ : Odrv12
    port map (
            O => \N__15749\,
            I => measured_delay_hc_11
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__15746\,
            I => measured_delay_hc_11
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__15737\,
            I => \N__15726\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__15736\,
            I => \N__15723\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__15735\,
            I => \N__15720\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__15734\,
            I => \N__15717\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__15733\,
            I => \N__15711\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__15732\,
            I => \N__15707\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__15731\,
            I => \N__15704\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15691\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15691\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15691\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15678\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15678\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15678\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15678\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15678\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15678\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15673\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15673\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15707\,
            I => \N__15666\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15666\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15666\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__15702\,
            I => \N__15662\
        );

    \I__3083\ : CascadeMux
    port map (
            O => \N__15701\,
            I => \N__15659\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__15700\,
            I => \N__15656\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__15699\,
            I => \N__15653\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15647\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15691\,
            I => \N__15644\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15678\,
            I => \N__15637\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15673\,
            I => \N__15637\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__15666\,
            I => \N__15637\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15634\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15618\
        );

    \I__3073\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15618\
        );

    \I__3072\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15618\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15618\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15618\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15618\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15618\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15615\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__15644\,
            I => \N__15608\
        );

    \I__3065\ : Span4Mux_v
    port map (
            O => \N__15637\,
            I => \N__15608\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15608\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15605\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__15618\,
            I => \N__15602\
        );

    \I__3061\ : Span4Mux_h
    port map (
            O => \N__15615\,
            I => \N__15599\
        );

    \I__3060\ : Span4Mux_h
    port map (
            O => \N__15608\,
            I => \N__15596\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__15605\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__3058\ : Odrv12
    port map (
            O => \N__15602\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__15599\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__15596\,
            I => \phase_controller_slave.start_timer_hcZ0\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15581\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15581\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15581\,
            I => \N__15573\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15566\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15566\
        );

    \I__3050\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15566\
        );

    \I__3049\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15563\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15576\,
            I => \N__15555\
        );

    \I__3047\ : Span4Mux_h
    port map (
            O => \N__15573\,
            I => \N__15548\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__15566\,
            I => \N__15548\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15563\,
            I => \N__15545\
        );

    \I__3044\ : InMux
    port map (
            O => \N__15562\,
            I => \N__15534\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15534\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15534\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15534\
        );

    \I__3040\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15534\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15527\
        );

    \I__3038\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15522\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15522\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__15548\,
            I => \N__15515\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__15545\,
            I => \N__15515\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__15534\,
            I => \N__15515\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15506\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15506\
        );

    \I__3031\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15506\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15506\
        );

    \I__3029\ : Odrv12
    port map (
            O => \N__15527\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15522\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__15515\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__15506\,
            I => \phase_controller_inst1.stoper_hc.un1_start\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15494\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__3023\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15488\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__15485\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__3020\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__15476\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__3017\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15470\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__15470\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15457\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15457\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15465\,
            I => \N__15440\
        );

    \I__3012\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15440\
        );

    \I__3011\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15440\
        );

    \I__3010\ : InMux
    port map (
            O => \N__15462\,
            I => \N__15440\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15457\,
            I => \N__15431\
        );

    \I__3008\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15420\
        );

    \I__3007\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15420\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15420\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15420\
        );

    \I__3004\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15420\
        );

    \I__3003\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15413\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15413\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15449\,
            I => \N__15413\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15408\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15395\
        );

    \I__2998\ : InMux
    port map (
            O => \N__15438\,
            I => \N__15395\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15437\,
            I => \N__15395\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15395\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15435\,
            I => \N__15395\
        );

    \I__2994\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15395\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__15431\,
            I => \N__15388\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__15420\,
            I => \N__15388\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__15413\,
            I => \N__15388\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15383\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15383\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__15408\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_d\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__15395\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_d\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__15388\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_d\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__15383\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_d\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \N__15370\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__15373\,
            I => \N__15367\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15362\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15362\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15362\,
            I => \N__15346\
        );

    \I__2979\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15337\
        );

    \I__2978\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15337\
        );

    \I__2977\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15337\
        );

    \I__2976\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15337\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__15357\,
            I => \N__15334\
        );

    \I__2974\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15318\
        );

    \I__2973\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15318\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15354\,
            I => \N__15318\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15318\
        );

    \I__2970\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15318\
        );

    \I__2969\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15311\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15311\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15311\
        );

    \I__2966\ : Span4Mux_v
    port map (
            O => \N__15346\,
            I => \N__15306\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__15337\,
            I => \N__15303\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15290\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15290\
        );

    \I__2962\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15290\
        );

    \I__2961\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15290\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15290\
        );

    \I__2959\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15290\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15285\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__15311\,
            I => \N__15285\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15280\
        );

    \I__2955\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15280\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__15306\,
            I => \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__15303\,
            I => \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__15290\,
            I => \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__15285\,
            I => \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__15280\,
            I => \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\
        );

    \I__2949\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15266\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__15266\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__15263\,
            I => \N__15251\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__15262\,
            I => \N__15248\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__15261\,
            I => \N__15245\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__15260\,
            I => \N__15242\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__15259\,
            I => \N__15239\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15258\,
            I => \N__15224\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15257\,
            I => \N__15215\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15215\
        );

    \I__2939\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15215\
        );

    \I__2938\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15215\
        );

    \I__2937\ : InMux
    port map (
            O => \N__15251\,
            I => \N__15212\
        );

    \I__2936\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15203\
        );

    \I__2935\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15203\
        );

    \I__2934\ : InMux
    port map (
            O => \N__15242\,
            I => \N__15203\
        );

    \I__2933\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15203\
        );

    \I__2932\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15200\
        );

    \I__2931\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15197\
        );

    \I__2930\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15190\
        );

    \I__2929\ : InMux
    port map (
            O => \N__15235\,
            I => \N__15190\
        );

    \I__2928\ : InMux
    port map (
            O => \N__15234\,
            I => \N__15190\
        );

    \I__2927\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15175\
        );

    \I__2926\ : InMux
    port map (
            O => \N__15232\,
            I => \N__15175\
        );

    \I__2925\ : InMux
    port map (
            O => \N__15231\,
            I => \N__15175\
        );

    \I__2924\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15175\
        );

    \I__2923\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15175\
        );

    \I__2922\ : InMux
    port map (
            O => \N__15228\,
            I => \N__15175\
        );

    \I__2921\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15175\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__15224\,
            I => \N__15172\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15165\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__15212\,
            I => \N__15165\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__15203\,
            I => \N__15158\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__15200\,
            I => \N__15158\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__15197\,
            I => \N__15158\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__15190\,
            I => \N__15153\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15153\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__15172\,
            I => \N__15150\
        );

    \I__2911\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15147\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15144\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__15165\,
            I => \N__15141\
        );

    \I__2908\ : Span12Mux_h
    port map (
            O => \N__15158\,
            I => \N__15138\
        );

    \I__2907\ : Span4Mux_v
    port map (
            O => \N__15153\,
            I => \N__15131\
        );

    \I__2906\ : Span4Mux_h
    port map (
            O => \N__15150\,
            I => \N__15131\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__15147\,
            I => \N__15131\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__15144\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__15141\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2902\ : Odrv12
    port map (
            O => \N__15138\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__15131\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\
        );

    \I__2900\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15119\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__15119\,
            I => \N__15115\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15112\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__15115\,
            I => \N__15106\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__15112\,
            I => \N__15106\
        );

    \I__2895\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15103\
        );

    \I__2894\ : Span4Mux_h
    port map (
            O => \N__15106\,
            I => \N__15098\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15095\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15090\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15090\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__15098\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__15095\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__15090\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__15083\,
            I => \N__15080\
        );

    \I__2886\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15058\
        );

    \I__2885\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15053\
        );

    \I__2884\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15053\
        );

    \I__2883\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15036\
        );

    \I__2882\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15036\
        );

    \I__2881\ : InMux
    port map (
            O => \N__15075\,
            I => \N__15036\
        );

    \I__2880\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15036\
        );

    \I__2879\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15036\
        );

    \I__2878\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15036\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15071\,
            I => \N__15036\
        );

    \I__2876\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15036\
        );

    \I__2875\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15033\
        );

    \I__2874\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15016\
        );

    \I__2873\ : InMux
    port map (
            O => \N__15067\,
            I => \N__15016\
        );

    \I__2872\ : InMux
    port map (
            O => \N__15066\,
            I => \N__15016\
        );

    \I__2871\ : InMux
    port map (
            O => \N__15065\,
            I => \N__15016\
        );

    \I__2870\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15016\
        );

    \I__2869\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15016\
        );

    \I__2868\ : InMux
    port map (
            O => \N__15062\,
            I => \N__15016\
        );

    \I__2867\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15016\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__15058\,
            I => \N__15009\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__15053\,
            I => \N__15009\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__15036\,
            I => \N__15009\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__15033\,
            I => \N__15003\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__15016\,
            I => \N__15003\
        );

    \I__2861\ : Span4Mux_v
    port map (
            O => \N__15009\,
            I => \N__14998\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__15008\,
            I => \N__14994\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__15003\,
            I => \N__14991\
        );

    \I__2858\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14988\
        );

    \I__2857\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14985\
        );

    \I__2856\ : Span4Mux_h
    port map (
            O => \N__14998\,
            I => \N__14982\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14979\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14976\
        );

    \I__2853\ : Sp12to4
    port map (
            O => \N__14991\,
            I => \N__14971\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14988\,
            I => \N__14971\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__14985\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__2850\ : Odrv4
    port map (
            O => \N__14982\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14979\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__14976\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__2847\ : Odrv12
    port map (
            O => \N__14971\,
            I => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14957\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__14957\,
            I => \N__14954\
        );

    \I__2844\ : Span4Mux_h
    port map (
            O => \N__14954\,
            I => \N__14950\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__14953\,
            I => \N__14947\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__14950\,
            I => \N__14942\
        );

    \I__2841\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14937\
        );

    \I__2840\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14937\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14934\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__14942\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14937\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__14934\,
            I => \phase_controller_slave.stoper_tr.time_passed11\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__14924\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__14921\,
            I => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14912\,
            I => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14906\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_0\
        );

    \I__2827\ : InMux
    port map (
            O => \N__14903\,
            I => \N__14897\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14902\,
            I => \N__14897\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14897\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14891\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__2822\ : Span4Mux_v
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__2821\ : Sp12to4
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__2820\ : Span12Mux_h
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__2819\ : Odrv12
    port map (
            O => \N__14879\,
            I => il_min_comp2_c
        );

    \I__2818\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14870\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14867\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14864\
        );

    \I__2815\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14860\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14870\,
            I => \N__14857\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14852\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__14864\,
            I => \N__14852\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14849\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14846\
        );

    \I__2809\ : Span4Mux_h
    port map (
            O => \N__14857\,
            I => \N__14843\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__14852\,
            I => \N__14840\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__14849\,
            I => measured_delay_hc_16
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__14846\,
            I => measured_delay_hc_16
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__14843\,
            I => measured_delay_hc_16
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__14840\,
            I => measured_delay_hc_16
        );

    \I__2803\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14825\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14821\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14818\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14815\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14811\
        );

    \I__2798\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14808\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__14821\,
            I => \N__14803\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__14818\,
            I => \N__14803\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14815\,
            I => \N__14800\
        );

    \I__2794\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14797\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__14811\,
            I => \N__14794\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__14808\,
            I => \N__14789\
        );

    \I__2791\ : Span4Mux_h
    port map (
            O => \N__14803\,
            I => \N__14789\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__14800\,
            I => \N__14786\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14797\,
            I => measured_delay_hc_14
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__14794\,
            I => measured_delay_hc_14
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__14789\,
            I => measured_delay_hc_14
        );

    \I__2786\ : Odrv4
    port map (
            O => \N__14786\,
            I => measured_delay_hc_14
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__14777\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__14771\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14768\,
            I => \N__14765\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14765\,
            I => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14756\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__14753\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_1\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__14747\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_\
        );

    \I__2773\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__14738\,
            I => \N__14735\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__14735\,
            I => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14726\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14723\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__14730\,
            I => \N__14719\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__14729\,
            I => \N__14716\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14711\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14711\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14708\
        );

    \I__2763\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14705\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14702\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__14711\,
            I => \N__14699\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__14708\,
            I => \N__14696\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__14705\,
            I => \N__14693\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__14702\,
            I => measured_delay_hc_5
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__14699\,
            I => measured_delay_hc_5
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__14696\,
            I => measured_delay_hc_5
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__14693\,
            I => measured_delay_hc_5
        );

    \I__2754\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14677\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14677\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14674\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14677\,
            I => \N__14671\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__14674\,
            I => measured_delay_hc_20
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__14671\,
            I => measured_delay_hc_20
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__14666\,
            I => \N__14662\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14659\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14656\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__14659\,
            I => \N__14653\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__14656\,
            I => \N__14647\
        );

    \I__2743\ : Span4Mux_h
    port map (
            O => \N__14653\,
            I => \N__14644\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14641\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14638\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14635\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__14647\,
            I => \N__14632\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__14644\,
            I => \N__14625\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14625\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14638\,
            I => \N__14625\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14635\,
            I => measured_delay_hc_3
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__14632\,
            I => measured_delay_hc_3
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__14625\,
            I => measured_delay_hc_3
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__14618\,
            I => \N__14611\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14608\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14605\
        );

    \I__2729\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14602\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14599\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14611\,
            I => \N__14596\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14608\,
            I => \N__14593\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__14605\,
            I => \N__14588\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14602\,
            I => \N__14588\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14599\,
            I => \N__14585\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14596\,
            I => \N__14580\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__14593\,
            I => \N__14580\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__14588\,
            I => \N__14577\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__14585\,
            I => measured_delay_hc_17
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__14580\,
            I => measured_delay_hc_17
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__14577\,
            I => measured_delay_hc_17
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__14570\,
            I => \N__14566\
        );

    \I__2715\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14562\
        );

    \I__2714\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14559\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14555\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__14562\,
            I => \N__14551\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__14559\,
            I => \N__14548\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__14558\,
            I => \N__14545\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__14555\,
            I => \N__14542\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14554\,
            I => \N__14539\
        );

    \I__2707\ : Span4Mux_v
    port map (
            O => \N__14551\,
            I => \N__14536\
        );

    \I__2706\ : Span4Mux_v
    port map (
            O => \N__14548\,
            I => \N__14533\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14530\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__14542\,
            I => \N__14525\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14539\,
            I => \N__14525\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__14536\,
            I => \N__14520\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__14533\,
            I => \N__14520\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__14530\,
            I => \N__14515\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__14525\,
            I => \N__14515\
        );

    \I__2698\ : Odrv4
    port map (
            O => \N__14520\,
            I => measured_delay_hc_6
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__14515\,
            I => measured_delay_hc_6
        );

    \I__2696\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14504\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14501\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__14508\,
            I => \N__14498\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14494\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14504\,
            I => \N__14489\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__14501\,
            I => \N__14489\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14486\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__14497\,
            I => \N__14483\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14494\,
            I => \N__14480\
        );

    \I__2687\ : Span4Mux_h
    port map (
            O => \N__14489\,
            I => \N__14475\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14475\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14472\
        );

    \I__2684\ : Span4Mux_h
    port map (
            O => \N__14480\,
            I => \N__14469\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__14475\,
            I => \N__14466\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__14472\,
            I => measured_delay_hc_13
        );

    \I__2681\ : Odrv4
    port map (
            O => \N__14469\,
            I => measured_delay_hc_13
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__14466\,
            I => measured_delay_hc_13
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__14459\,
            I => \N__14454\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__14458\,
            I => \N__14451\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14446\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14443\
        );

    \I__2675\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14440\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__14450\,
            I => \N__14437\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14434\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__14446\,
            I => \N__14431\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__14443\,
            I => \N__14428\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__14440\,
            I => \N__14425\
        );

    \I__2669\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14422\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__14434\,
            I => \N__14419\
        );

    \I__2667\ : Span4Mux_v
    port map (
            O => \N__14431\,
            I => \N__14416\
        );

    \I__2666\ : Span4Mux_h
    port map (
            O => \N__14428\,
            I => \N__14413\
        );

    \I__2665\ : Span4Mux_v
    port map (
            O => \N__14425\,
            I => \N__14410\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__14422\,
            I => measured_delay_hc_19
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__14419\,
            I => measured_delay_hc_19
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__14416\,
            I => measured_delay_hc_19
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__14413\,
            I => measured_delay_hc_19
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__14410\,
            I => measured_delay_hc_19
        );

    \I__2659\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14394\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14389\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__14397\,
            I => \N__14386\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__14394\,
            I => \N__14382\
        );

    \I__2655\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14379\
        );

    \I__2654\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14376\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14373\
        );

    \I__2652\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14370\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__14385\,
            I => \N__14367\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__14382\,
            I => \N__14360\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__14379\,
            I => \N__14360\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__14376\,
            I => \N__14360\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__14373\,
            I => \N__14355\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__14370\,
            I => \N__14355\
        );

    \I__2645\ : InMux
    port map (
            O => \N__14367\,
            I => \N__14352\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__14360\,
            I => \N__14349\
        );

    \I__2643\ : Span4Mux_h
    port map (
            O => \N__14355\,
            I => \N__14346\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__14352\,
            I => measured_delay_hc_15
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__14349\,
            I => measured_delay_hc_15
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__14346\,
            I => measured_delay_hc_15
        );

    \I__2639\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14334\
        );

    \I__2638\ : InMux
    port map (
            O => \N__14338\,
            I => \N__14329\
        );

    \I__2637\ : InMux
    port map (
            O => \N__14337\,
            I => \N__14326\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14334\,
            I => \N__14323\
        );

    \I__2635\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14320\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14332\,
            I => \N__14317\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14329\,
            I => \N__14308\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__14326\,
            I => \N__14308\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__14323\,
            I => \N__14308\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__14320\,
            I => \N__14308\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14317\,
            I => \N__14305\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__14308\,
            I => \N__14302\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__14305\,
            I => measured_delay_hc_18
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__14302\,
            I => measured_delay_hc_18
        );

    \I__2625\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14294\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14294\,
            I => \N__14291\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__14291\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__14285\,
            I => \N__14282\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__14282\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14276\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__14273\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__2616\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14267\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__14267\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14264\,
            I => \N__14259\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14256\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14253\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__14259\,
            I => \N__14246\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__14256\,
            I => \N__14246\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14253\,
            I => \N__14243\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14240\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14237\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__14246\,
            I => \N__14234\
        );

    \I__2605\ : Span4Mux_h
    port map (
            O => \N__14243\,
            I => \N__14229\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__14240\,
            I => \N__14229\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__14237\,
            I => measured_delay_hc_4
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__14234\,
            I => measured_delay_hc_4
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__14229\,
            I => measured_delay_hc_4
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__14222\,
            I => \N__14218\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__14221\,
            I => \N__14215\
        );

    \I__2598\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14211\
        );

    \I__2597\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14208\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__14214\,
            I => \N__14203\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__14211\,
            I => \N__14200\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__14208\,
            I => \N__14197\
        );

    \I__2593\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14192\
        );

    \I__2592\ : InMux
    port map (
            O => \N__14206\,
            I => \N__14192\
        );

    \I__2591\ : InMux
    port map (
            O => \N__14203\,
            I => \N__14189\
        );

    \I__2590\ : Span4Mux_h
    port map (
            O => \N__14200\,
            I => \N__14186\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__14197\,
            I => \N__14183\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14180\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__14189\,
            I => measured_delay_hc_1
        );

    \I__2586\ : Odrv4
    port map (
            O => \N__14186\,
            I => measured_delay_hc_1
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__14183\,
            I => measured_delay_hc_1
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__14180\,
            I => measured_delay_hc_1
        );

    \I__2583\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14164\
        );

    \I__2582\ : InMux
    port map (
            O => \N__14170\,
            I => \N__14164\
        );

    \I__2581\ : InMux
    port map (
            O => \N__14169\,
            I => \N__14161\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14153\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__14158\,
            I => \N__14153\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__14153\,
            I => measured_delay_hc_22
        );

    \I__2576\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14143\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14143\
        );

    \I__2574\ : InMux
    port map (
            O => \N__14148\,
            I => \N__14140\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__14143\,
            I => \N__14137\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__14140\,
            I => \N__14132\
        );

    \I__2571\ : Span4Mux_h
    port map (
            O => \N__14137\,
            I => \N__14132\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__14132\,
            I => measured_delay_hc_21
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__14129\,
            I => \N__14126\
        );

    \I__2568\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14123\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__14123\,
            I => \N__14117\
        );

    \I__2566\ : InMux
    port map (
            O => \N__14122\,
            I => \N__14114\
        );

    \I__2565\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14111\
        );

    \I__2564\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14108\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__14117\,
            I => \N__14105\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__14114\,
            I => \N__14102\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__14111\,
            I => \N__14099\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__14108\,
            I => measured_delay_hc_0
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__14105\,
            I => measured_delay_hc_0
        );

    \I__2558\ : Odrv12
    port map (
            O => \N__14102\,
            I => measured_delay_hc_0
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__14099\,
            I => measured_delay_hc_0
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__2555\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14084\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__14084\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__14081\,
            I => \N__14078\
        );

    \I__2552\ : InMux
    port map (
            O => \N__14078\,
            I => \N__14075\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__14075\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__14072\,
            I => \N__14069\
        );

    \I__2549\ : InMux
    port map (
            O => \N__14069\,
            I => \N__14066\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__14066\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\
        );

    \I__2547\ : CascadeMux
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__2546\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14057\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__14057\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\
        );

    \I__2544\ : InMux
    port map (
            O => \N__14054\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__14051\,
            I => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\
        );

    \I__2542\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14045\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__14045\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__14042\,
            I => \N__14039\
        );

    \I__2539\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14036\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__14036\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__14033\,
            I => \N__14030\
        );

    \I__2536\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14027\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__14027\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2533\ : InMux
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__14018\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__2530\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__14009\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__2527\ : InMux
    port map (
            O => \N__14003\,
            I => \N__14000\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__14000\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13994\,
            I => \N__13991\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__13991\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13982\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13973\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__13973\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__13967\,
            I => \N__13964\
        );

    \I__2514\ : Span4Mux_h
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__13961\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__13958\,
            I => \N__13955\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__13952\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__13949\,
            I => \N__13946\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13943\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__13943\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\
        );

    \I__2506\ : InMux
    port map (
            O => \N__13940\,
            I => \N__13937\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13937\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__13934\,
            I => \N__13931\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13928\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__13928\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13922\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13922\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13916\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13913\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__13913\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13910\,
            I => \N__13907\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13907\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13898\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13898\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__13889\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__2487\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__13880\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13874\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__13871\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13862\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__13853\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__13850\,
            I => \N__13847\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__13844\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__13835\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__13832\,
            I => \N__13829\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13826\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__2467\ : CEMux
    port map (
            O => \N__13823\,
            I => \N__13819\
        );

    \I__2466\ : CEMux
    port map (
            O => \N__13822\,
            I => \N__13816\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13819\,
            I => \N__13813\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__13816\,
            I => \N__13809\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__13813\,
            I => \N__13806\
        );

    \I__2462\ : CEMux
    port map (
            O => \N__13812\,
            I => \N__13803\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__13809\,
            I => \N__13800\
        );

    \I__2460\ : Span4Mux_s2_h
    port map (
            O => \N__13806\,
            I => \N__13795\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13803\,
            I => \N__13795\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__13800\,
            I => \N__13792\
        );

    \I__2457\ : Sp12to4
    port map (
            O => \N__13795\,
            I => \N__13789\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__13792\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__13789\,
            I => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__13784\,
            I => \N__13779\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13776\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13773\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13770\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__13776\,
            I => \N__13766\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13773\,
            I => \N__13763\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13770\,
            I => \N__13760\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__13769\,
            I => \N__13757\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__13766\,
            I => \N__13754\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__13763\,
            I => \N__13749\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__13760\,
            I => \N__13749\
        );

    \I__2443\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13746\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__13754\,
            I => measured_delay_tr_19
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__13749\,
            I => measured_delay_tr_19
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13746\,
            I => measured_delay_tr_19
        );

    \I__2439\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13736\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__13736\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13729\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__13729\,
            I => \N__13723\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13726\,
            I => \N__13720\
        );

    \I__2433\ : Span4Mux_h
    port map (
            O => \N__13723\,
            I => \N__13715\
        );

    \I__2432\ : Span4Mux_h
    port map (
            O => \N__13720\,
            I => \N__13712\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13709\
        );

    \I__2430\ : InMux
    port map (
            O => \N__13718\,
            I => \N__13706\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__13715\,
            I => measured_delay_tr_17
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__13712\,
            I => measured_delay_tr_17
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__13709\,
            I => measured_delay_tr_17
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__13706\,
            I => measured_delay_tr_17
        );

    \I__2425\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13694\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13694\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13687\
        );

    \I__2422\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13684\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__13687\,
            I => \N__13681\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__13684\,
            I => \N__13678\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__13681\,
            I => \N__13671\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__13678\,
            I => \N__13671\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13668\
        );

    \I__2416\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13665\
        );

    \I__2415\ : Odrv4
    port map (
            O => \N__13671\,
            I => measured_delay_tr_18
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__13668\,
            I => measured_delay_tr_18
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__13665\,
            I => measured_delay_tr_18
        );

    \I__2412\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13655\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N__13645\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13648\,
            I => \N__13641\
        );

    \I__2407\ : Span4Mux_h
    port map (
            O => \N__13645\,
            I => \N__13637\
        );

    \I__2406\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13634\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__13641\,
            I => \N__13631\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13628\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__13637\,
            I => \N__13623\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__13634\,
            I => \N__13623\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__13631\,
            I => measured_delay_tr_16
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__13628\,
            I => measured_delay_tr_16
        );

    \I__2399\ : Odrv4
    port map (
            O => \N__13623\,
            I => measured_delay_tr_16
        );

    \I__2398\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__2396\ : Odrv12
    port map (
            O => \N__13610\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13595\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13595\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13595\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13595\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__2390\ : Span4Mux_h
    port map (
            O => \N__13592\,
            I => \N__13585\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13591\,
            I => \N__13576\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13576\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13576\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13576\
        );

    \I__2385\ : Span4Mux_v
    port map (
            O => \N__13585\,
            I => \N__13573\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__13576\,
            I => \N__13570\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__13573\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__2382\ : Odrv12
    port map (
            O => \N__13570\,
            I => \phase_controller_inst1.stoper_hc.un2_startlt31\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__13565\,
            I => \N__13562\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13559\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13556\,
            I => \N__13553\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__13550\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13541\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__13538\,
            I => \N__13535\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13532\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13532\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__13529\,
            I => \N__13526\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13526\,
            I => \N__13523\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13523\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__2365\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13514\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__13511\,
            I => \N__13508\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__13505\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__13502\,
            I => \N__13499\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13496\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__13496\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13493\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__13484\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__13481\,
            I => \N__13478\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__13475\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__13469\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13460\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13460\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__13451\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__2341\ : InMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__13442\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__13433\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__13424\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13421\,
            I => \N__13418\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__13415\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__2329\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13406\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13406\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13400\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__13397\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__13394\,
            I => \N__13391\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13391\,
            I => \N__13388\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13388\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__2319\ : Odrv12
    port map (
            O => \N__13379\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2317\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13370\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__13370\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__2315\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13364\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__13361\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13355\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13355\,
            I => \N__13350\
        );

    \I__2310\ : InMux
    port map (
            O => \N__13354\,
            I => \N__13347\
        );

    \I__2309\ : InMux
    port map (
            O => \N__13353\,
            I => \N__13344\
        );

    \I__2308\ : Odrv12
    port map (
            O => \N__13350\,
            I => measured_delay_tr_2
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__13347\,
            I => measured_delay_tr_2
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__13344\,
            I => measured_delay_tr_2
        );

    \I__2305\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13331\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13331\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__13328\,
            I => \N__13322\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13317\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13317\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13325\,
            I => \N__13314\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__13322\,
            I => measured_delay_tr_3
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__13317\,
            I => measured_delay_tr_3
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13314\,
            I => measured_delay_tr_3
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__13307\,
            I => \N__13303\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13294\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13294\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13294\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__13301\,
            I => \N__13290\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13294\,
            I => \N__13286\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13279\
        );

    \I__2288\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13279\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13279\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__13286\,
            I => \N__13276\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__13279\,
            I => \N__13273\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__13276\,
            I => \phase_controller_inst1.stoper_tr.N_109\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__13273\,
            I => \phase_controller_inst1.stoper_tr.N_109\
        );

    \I__2282\ : InMux
    port map (
            O => \N__13268\,
            I => \N__13256\
        );

    \I__2281\ : InMux
    port map (
            O => \N__13267\,
            I => \N__13256\
        );

    \I__2280\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13256\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13249\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13249\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13249\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13246\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__13249\,
            I => \N__13243\
        );

    \I__2274\ : Span4Mux_h
    port map (
            O => \N__13246\,
            I => \N__13240\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__13243\,
            I => \phase_controller_inst1.stoper_tr.N_110\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__13240\,
            I => \phase_controller_inst1.stoper_tr.N_110\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__13235\,
            I => \N__13228\
        );

    \I__2270\ : CascadeMux
    port map (
            O => \N__13234\,
            I => \N__13225\
        );

    \I__2269\ : CascadeMux
    port map (
            O => \N__13233\,
            I => \N__13221\
        );

    \I__2268\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13218\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13231\,
            I => \N__13213\
        );

    \I__2266\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13213\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13208\
        );

    \I__2264\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13208\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13205\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__13218\,
            I => \N__13200\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__13213\,
            I => \N__13200\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__13208\,
            I => \N__13195\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__13205\,
            I => \N__13195\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__13200\,
            I => \N__13192\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__13195\,
            I => \phase_controller_inst1.stoper_tr.N_92\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__13192\,
            I => \phase_controller_inst1.stoper_tr.N_92\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \N__13184\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13180\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__13183\,
            I => \N__13176\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__13180\,
            I => \N__13173\
        );

    \I__2251\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13170\
        );

    \I__2250\ : InMux
    port map (
            O => \N__13176\,
            I => \N__13167\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__13173\,
            I => \N__13162\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__13170\,
            I => \N__13162\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__13167\,
            I => measured_delay_tr_6
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__13162\,
            I => measured_delay_tr_6
        );

    \I__2245\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13146\
        );

    \I__2244\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13146\
        );

    \I__2243\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13146\
        );

    \I__2242\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13141\
        );

    \I__2241\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13141\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__13146\,
            I => \N__13133\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__13141\,
            I => \N__13130\
        );

    \I__2238\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13119\
        );

    \I__2237\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13119\
        );

    \I__2236\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13119\
        );

    \I__2235\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13119\
        );

    \I__2234\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13119\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__13133\,
            I => \N__13115\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__13130\,
            I => \N__13110\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__13119\,
            I => \N__13110\
        );

    \I__2230\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13107\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__13115\,
            I => \phase_controller_inst1.stoper_tr.N_95\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__13110\,
            I => \phase_controller_inst1.stoper_tr.N_95\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__13107\,
            I => \phase_controller_inst1.stoper_tr.N_95\
        );

    \I__2226\ : InMux
    port map (
            O => \N__13100\,
            I => \N__13097\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__13097\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__13094\,
            I => \N__13091\
        );

    \I__2223\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13088\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__13088\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13082\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__13082\,
            I => \N__13079\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__13079\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__2217\ : InMux
    port map (
            O => \N__13073\,
            I => \N__13070\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__13070\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__2215\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__13064\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__13061\,
            I => \N__13058\
        );

    \I__2212\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13055\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__13055\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__2210\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13049\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__13049\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__13046\,
            I => \N__13043\
        );

    \I__2207\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13040\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__13040\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13037\,
            I => \N__13034\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__13034\,
            I => \N__13031\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__13031\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__13028\,
            I => \N__13025\
        );

    \I__2201\ : InMux
    port map (
            O => \N__13025\,
            I => \N__13022\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__13022\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__2199\ : InMux
    port map (
            O => \N__13019\,
            I => \N__13016\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__13016\,
            I => \N__13012\
        );

    \I__2197\ : InMux
    port map (
            O => \N__13015\,
            I => \N__13009\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__13012\,
            I => \N__13003\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__13009\,
            I => \N__13003\
        );

    \I__2194\ : InMux
    port map (
            O => \N__13008\,
            I => \N__13000\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__13003\,
            I => measured_delay_tr_12
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__13000\,
            I => measured_delay_tr_12
        );

    \I__2191\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12991\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12988\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12991\,
            I => \N__12984\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__12988\,
            I => \N__12981\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__12987\,
            I => \N__12978\
        );

    \I__2186\ : Span4Mux_h
    port map (
            O => \N__12984\,
            I => \N__12975\
        );

    \I__2185\ : Span4Mux_h
    port map (
            O => \N__12981\,
            I => \N__12972\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12969\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__12975\,
            I => measured_delay_tr_13
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__12972\,
            I => measured_delay_tr_13
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12969\,
            I => measured_delay_tr_13
        );

    \I__2180\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12958\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12953\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__12958\,
            I => \N__12949\
        );

    \I__2177\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12944\
        );

    \I__2176\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12944\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12953\,
            I => \N__12941\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12938\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__12949\,
            I => \N__12933\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12944\,
            I => \N__12933\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__12941\,
            I => measured_delay_tr_14
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12938\,
            I => measured_delay_tr_14
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__12933\,
            I => measured_delay_tr_14
        );

    \I__2168\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12911\
        );

    \I__2167\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12911\
        );

    \I__2166\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12911\
        );

    \I__2165\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12911\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12911\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12907\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__12910\,
            I => \N__12900\
        );

    \I__2161\ : Span4Mux_v
    port map (
            O => \N__12907\,
            I => \N__12897\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12906\,
            I => \N__12886\
        );

    \I__2159\ : InMux
    port map (
            O => \N__12905\,
            I => \N__12886\
        );

    \I__2158\ : InMux
    port map (
            O => \N__12904\,
            I => \N__12886\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12903\,
            I => \N__12886\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12900\,
            I => \N__12886\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__12897\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__12886\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12877\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12874\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__12877\,
            I => \N__12870\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12874\,
            I => \N__12867\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12864\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__12870\,
            I => measured_delay_tr_10
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__12867\,
            I => measured_delay_tr_10
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12864\,
            I => measured_delay_tr_10
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__12857\,
            I => \N__12853\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12850\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12847\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__12850\,
            I => \N__12844\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12840\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__12844\,
            I => \N__12837\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12843\,
            I => \N__12834\
        );

    \I__2138\ : Odrv12
    port map (
            O => \N__12840\,
            I => measured_delay_tr_4
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__12837\,
            I => measured_delay_tr_4
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12834\,
            I => measured_delay_tr_4
        );

    \I__2135\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12824\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__12824\,
            I => \N__12819\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12812\
        );

    \I__2132\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12812\
        );

    \I__2131\ : Span4Mux_v
    port map (
            O => \N__12819\,
            I => \N__12809\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12806\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__12817\,
            I => \N__12803\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__12812\,
            I => \N__12800\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__12809\,
            I => \N__12795\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12806\,
            I => \N__12795\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12792\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__12800\,
            I => \N__12789\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__12795\,
            I => measured_delay_tr_7
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__12792\,
            I => measured_delay_tr_7
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__12789\,
            I => measured_delay_tr_7
        );

    \I__2120\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12779\,
            I => \N__12773\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12778\,
            I => \N__12770\
        );

    \I__2117\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12767\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12776\,
            I => \N__12764\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__12773\,
            I => \N__12759\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__12770\,
            I => \N__12759\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__12767\,
            I => \N__12756\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12753\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__12759\,
            I => \N__12750\
        );

    \I__2110\ : Odrv12
    port map (
            O => \N__12756\,
            I => measured_delay_tr_8
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12753\,
            I => measured_delay_tr_8
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__12750\,
            I => measured_delay_tr_8
        );

    \I__2107\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__12740\,
            I => \N__12735\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12732\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12729\
        );

    \I__2103\ : Span4Mux_h
    port map (
            O => \N__12735\,
            I => \N__12724\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__12732\,
            I => \N__12724\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12729\,
            I => measured_delay_tr_5
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__12724\,
            I => measured_delay_tr_5
        );

    \I__2099\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12716\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__12713\,
            I => \N__12709\
        );

    \I__2096\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12706\
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__12709\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__12706\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__12701\,
            I => \N__12697\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__12700\,
            I => \N__12694\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12691\
        );

    \I__2090\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12688\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__12691\,
            I => \N__12685\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12688\,
            I => measured_delay_tr_1
        );

    \I__2087\ : Odrv12
    port map (
            O => \N__12685\,
            I => measured_delay_tr_1
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__12680\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3_cascade_\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12674\,
            I => \phase_controller_inst1.stoper_hc.un1_m2_eZ0\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__12671\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__12665\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__12662\,
            I => \N__12659\
        );

    \I__2079\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__12656\,
            I => \N__12652\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12649\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__12652\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__12649\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0\
        );

    \I__2074\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__12641\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12635\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__2070\ : Glb2LocalMux
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__2069\ : GlobalMux
    port map (
            O => \N__12629\,
            I => clk_12mhz
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__12626\,
            I => \N__12623\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12623\,
            I => \N__12620\
        );

    \I__2066\ : IoSpan4Mux
    port map (
            O => \N__12620\,
            I => \N__12617\
        );

    \I__2065\ : Span4Mux_s0_v
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__12614\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12607\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12604\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__12607\,
            I => \N__12600\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__12604\,
            I => \N__12597\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__12600\,
            I => measured_delay_tr_11
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__12597\,
            I => measured_delay_tr_11
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12594\,
            I => measured_delay_tr_11
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__12587\,
            I => \N__12583\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__12586\,
            I => \N__12580\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12583\,
            I => \N__12577\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12574\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12577\,
            I => \N__12571\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__12574\,
            I => \N__12568\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__12571\,
            I => \N__12563\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__12568\,
            I => \N__12560\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12567\,
            I => \N__12555\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12555\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__12563\,
            I => measured_delay_tr_9
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__12560\,
            I => measured_delay_tr_9
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12555\,
            I => measured_delay_tr_9
        );

    \I__2042\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12545\,
            I => \N__12541\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12538\
        );

    \I__2039\ : Span4Mux_h
    port map (
            O => \N__12541\,
            I => \N__12532\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12538\,
            I => \N__12529\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12522\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12522\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12522\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__12532\,
            I => \phase_controller_inst1.stoper_tr.N_98\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__12529\,
            I => \phase_controller_inst1.stoper_tr.N_98\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__12522\,
            I => \phase_controller_inst1.stoper_tr.N_98\
        );

    \I__2031\ : InMux
    port map (
            O => \N__12515\,
            I => \N__12511\
        );

    \I__2030\ : InMux
    port map (
            O => \N__12514\,
            I => \N__12508\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12511\,
            I => phase_controller_inst1_stoper_hc_un1_startlto19_2
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__12508\,
            I => phase_controller_inst1_stoper_hc_un1_startlto19_2
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \phase_controller_inst1_stoper_hc_un1_startlto19_2_cascade_\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__12500\,
            I => \N__12492\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__12499\,
            I => \N__12489\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__12498\,
            I => \N__12486\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__12497\,
            I => \N__12476\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__12496\,
            I => \N__12473\
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__12495\,
            I => \N__12470\
        );

    \I__2020\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12457\
        );

    \I__2019\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12457\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12457\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12448\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12448\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12483\,
            I => \N__12448\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12448\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12441\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12441\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12441\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12434\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12434\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12434\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12427\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12427\
        );

    \I__2005\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12427\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12424\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12421\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__12464\,
            I => \N__12418\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12457\,
            I => \N__12407\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12448\,
            I => \N__12407\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__12441\,
            I => \N__12407\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12434\,
            I => \N__12400\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12427\,
            I => \N__12400\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12424\,
            I => \N__12400\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12421\,
            I => \N__12397\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12418\,
            I => \N__12393\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12417\,
            I => \N__12388\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12388\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12383\
        );

    \I__1990\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12383\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__12407\,
            I => \N__12378\
        );

    \I__1988\ : Span4Mux_h
    port map (
            O => \N__12400\,
            I => \N__12378\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__12397\,
            I => \N__12375\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12372\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__12393\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__12388\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12383\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__12378\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__12375\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12372\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12326\
        );

    \I__1978\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12326\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12326\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12326\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12326\
        );

    \I__1974\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12326\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12326\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12319\
        );

    \I__1971\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12319\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12319\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12306\
        );

    \I__1968\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12306\
        );

    \I__1967\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12306\
        );

    \I__1966\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12306\
        );

    \I__1965\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12306\
        );

    \I__1964\ : InMux
    port map (
            O => \N__12344\,
            I => \N__12306\
        );

    \I__1963\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12303\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12300\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__12341\,
            I => \N__12297\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__12326\,
            I => \N__12288\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__12319\,
            I => \N__12288\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12283\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12283\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__12300\,
            I => \N__12280\
        );

    \I__1955\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12274\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12296\,
            I => \N__12274\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12267\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12267\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12267\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__12288\,
            I => \N__12262\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__12283\,
            I => \N__12262\
        );

    \I__1948\ : Span4Mux_h
    port map (
            O => \N__12280\,
            I => \N__12259\
        );

    \I__1947\ : InMux
    port map (
            O => \N__12279\,
            I => \N__12256\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12274\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__12267\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__12262\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__12259\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__12256\,
            I => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\
        );

    \I__1941\ : CEMux
    port map (
            O => \N__12245\,
            I => \N__12242\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__12242\,
            I => \N__12236\
        );

    \I__1939\ : CEMux
    port map (
            O => \N__12241\,
            I => \N__12233\
        );

    \I__1938\ : CEMux
    port map (
            O => \N__12240\,
            I => \N__12230\
        );

    \I__1937\ : CEMux
    port map (
            O => \N__12239\,
            I => \N__12227\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__12236\,
            I => \N__12224\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__12233\,
            I => \N__12221\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12218\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__12227\,
            I => \N__12215\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__12224\,
            I => \N__12212\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__12221\,
            I => \N__12209\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__12218\,
            I => \N__12206\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__12215\,
            I => \N__12203\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__12212\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__12209\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__12206\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__12203\,
            I => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\
        );

    \I__1924\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__12191\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_a0Z0Z_1\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__12188\,
            I => \phase_controller_inst1.stoper_hc.un1_startlto31_aZ0Z2_cascade_\
        );

    \I__1921\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12181\
        );

    \I__1920\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__12181\,
            I => \d_N_5_mux\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__12178\,
            I => \d_N_5_mux\
        );

    \I__1917\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12170\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__12167\,
            I => \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__12164\,
            I => \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_2_cascade_\
        );

    \I__1913\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12157\
        );

    \I__1912\ : InMux
    port map (
            O => \N__12160\,
            I => \N__12154\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__12157\,
            I => \N__12151\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__12154\,
            I => \phase_controller_inst1.stoper_hc.un1_N_6_mux\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__12151\,
            I => \phase_controller_inst1.stoper_hc.un1_N_6_mux\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__12146\,
            I => \N__12143\
        );

    \I__1907\ : InMux
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__12140\,
            I => \phase_controller_inst1.stoper_hc.un1_m3_eZ0Z_1\
        );

    \I__1905\ : InMux
    port map (
            O => \N__12137\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__12134\,
            I => \N__12129\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__12133\,
            I => \N__12126\
        );

    \I__1902\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12123\
        );

    \I__1901\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12118\
        );

    \I__1900\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12118\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__12123\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__12118\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__1897\ : InMux
    port map (
            O => \N__12113\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__12110\,
            I => \N__12105\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__12109\,
            I => \N__12102\
        );

    \I__1894\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12099\
        );

    \I__1893\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12094\
        );

    \I__1892\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12094\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__12099\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__12094\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__1889\ : InMux
    port map (
            O => \N__12089\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__1888\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12081\
        );

    \I__1887\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12078\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12075\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__12081\,
            I => \N__12072\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__12078\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__12075\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__12072\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__1881\ : InMux
    port map (
            O => \N__12065\,
            I => \bfn_5_18_0_\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12057\
        );

    \I__1879\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12054\
        );

    \I__1878\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12051\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__12057\,
            I => \N__12048\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__12054\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__12051\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__12048\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__1873\ : InMux
    port map (
            O => \N__12041\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__12038\,
            I => \N__12033\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__12037\,
            I => \N__12030\
        );

    \I__1870\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12027\
        );

    \I__1869\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12022\
        );

    \I__1868\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12022\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__12027\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__12022\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__1865\ : InMux
    port map (
            O => \N__12017\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__12014\,
            I => \N__12009\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__12013\,
            I => \N__12006\
        );

    \I__1862\ : InMux
    port map (
            O => \N__12012\,
            I => \N__12003\
        );

    \I__1861\ : InMux
    port map (
            O => \N__12009\,
            I => \N__11998\
        );

    \I__1860\ : InMux
    port map (
            O => \N__12006\,
            I => \N__11998\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__12003\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11998\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11993\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11986\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11983\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__11986\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__11983\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11978\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11937\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11937\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11973\,
            I => \N__11937\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11937\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11971\,
            I => \N__11928\
        );

    \I__1846\ : InMux
    port map (
            O => \N__11970\,
            I => \N__11928\
        );

    \I__1845\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11928\
        );

    \I__1844\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11928\
        );

    \I__1843\ : InMux
    port map (
            O => \N__11967\,
            I => \N__11923\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11966\,
            I => \N__11923\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11965\,
            I => \N__11914\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11914\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11914\
        );

    \I__1838\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11914\
        );

    \I__1837\ : InMux
    port map (
            O => \N__11961\,
            I => \N__11905\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11905\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11905\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11905\
        );

    \I__1833\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11896\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11896\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11896\
        );

    \I__1830\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11896\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11887\
        );

    \I__1828\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11887\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11887\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11950\,
            I => \N__11887\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11949\,
            I => \N__11878\
        );

    \I__1824\ : InMux
    port map (
            O => \N__11948\,
            I => \N__11878\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11878\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11946\,
            I => \N__11878\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11937\,
            I => \N__11875\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11928\,
            I => \N__11860\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11923\,
            I => \N__11860\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11914\,
            I => \N__11860\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11860\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11896\,
            I => \N__11860\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__11887\,
            I => \N__11860\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11860\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__11875\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__1812\ : Odrv12
    port map (
            O => \N__11860\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11855\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11848\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11845\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11848\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__11845\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__1806\ : CEMux
    port map (
            O => \N__11840\,
            I => \N__11828\
        );

    \I__1805\ : CEMux
    port map (
            O => \N__11839\,
            I => \N__11828\
        );

    \I__1804\ : CEMux
    port map (
            O => \N__11838\,
            I => \N__11828\
        );

    \I__1803\ : CEMux
    port map (
            O => \N__11837\,
            I => \N__11828\
        );

    \I__1802\ : GlobalMux
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__1801\ : gio2CtrlBuf
    port map (
            O => \N__11825\,
            I => \delay_measurement_inst.delay_tr_timer.N_139_i_g\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11817\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11812\
        );

    \I__1798\ : InMux
    port map (
            O => \N__11820\,
            I => \N__11812\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__11817\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__11812\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11807\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__11804\,
            I => \N__11799\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__11803\,
            I => \N__11796\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11793\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11788\
        );

    \I__1790\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11788\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__11793\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__11788\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11783\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11780\,
            I => \N__11775\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \N__11772\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11769\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11764\
        );

    \I__1782\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11764\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__11769\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11764\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11759\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11751\
        );

    \I__1777\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11748\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11745\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11742\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11748\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__11745\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__11742\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11735\,
            I => \bfn_5_17_0_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11727\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11724\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11721\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11727\,
            I => \N__11718\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11724\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__11721\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__11718\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11711\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__11708\,
            I => \N__11703\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__11707\,
            I => \N__11700\
        );

    \I__1760\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11697\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11692\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11692\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__11697\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__11692\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11687\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__11684\,
            I => \N__11679\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__11683\,
            I => \N__11676\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11682\,
            I => \N__11673\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11668\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11668\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11673\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__11668\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__1747\ : InMux
    port map (
            O => \N__11663\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11655\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11650\
        );

    \I__1744\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11650\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__11655\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__11650\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__1741\ : InMux
    port map (
            O => \N__11645\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__1740\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11637\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11632\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11640\,
            I => \N__11632\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__11637\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11632\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11622\
        );

    \I__1734\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11617\
        );

    \I__1733\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11617\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__11622\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__11617\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11612\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__11609\,
            I => \N__11604\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \N__11601\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11598\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11593\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11593\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__11598\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__11593\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11588\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__11585\,
            I => \N__11580\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11584\,
            I => \N__11577\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11574\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11569\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11577\,
            I => \N__11569\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11574\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11569\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11564\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__1713\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11556\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11553\
        );

    \I__1711\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11550\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__11556\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__11553\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11550\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__1707\ : InMux
    port map (
            O => \N__11543\,
            I => \bfn_5_16_0_\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11535\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11532\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11529\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11535\,
            I => \N__11526\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11532\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__11529\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__11526\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__1699\ : InMux
    port map (
            O => \N__11519\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__11516\,
            I => \N__11511\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__11515\,
            I => \N__11508\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11505\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11500\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11500\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11505\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__11500\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__1691\ : InMux
    port map (
            O => \N__11495\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__11492\,
            I => \N__11487\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__11491\,
            I => \N__11484\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11481\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11476\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11476\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__11481\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11476\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__1683\ : InMux
    port map (
            O => \N__11471\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11468\,
            I => \N__11463\
        );

    \I__1681\ : InMux
    port map (
            O => \N__11467\,
            I => \N__11458\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11458\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__11463\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11458\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11453\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11450\,
            I => \N__11445\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11440\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11440\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11445\,
            I => \N__11437\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11434\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__11437\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__11434\,
            I => \delay_measurement_inst.elapsed_time_tr_18\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__11429\,
            I => \N__11424\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11421\
        );

    \I__1667\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11416\
        );

    \I__1666\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11416\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__11421\,
            I => \N__11413\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11410\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__11413\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__11410\,
            I => \delay_measurement_inst.elapsed_time_tr_19\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__11405\,
            I => \N__11401\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11397\
        );

    \I__1659\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11392\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11392\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__11397\,
            I => \N__11389\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__11392\,
            I => \N__11386\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__11389\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__11386\,
            I => \delay_measurement_inst.elapsed_time_tr_17\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11370\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11370\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11370\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11365\
        );

    \I__1649\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11365\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11370\,
            I => \N__11357\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__11365\,
            I => \N__11354\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11347\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11347\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11347\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11342\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11342\
        );

    \I__1641\ : Span4Mux_h
    port map (
            O => \N__11357\,
            I => \N__11339\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__11354\,
            I => \N__11336\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11347\,
            I => \N__11331\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11331\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__11339\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__11336\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__1635\ : Odrv12
    port map (
            O => \N__11331\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\
        );

    \I__1634\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11315\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11315\
        );

    \I__1632\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11308\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11308\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11308\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__11315\,
            I => \delay_measurement_inst.N_197_1\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__11308\,
            I => \delay_measurement_inst.N_197_1\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__11303\,
            I => \N__11299\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11296\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__11290\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__1621\ : Odrv4
    port map (
            O => \N__11287\,
            I => \delay_measurement_inst.elapsed_time_tr_13\
        );

    \I__1620\ : CEMux
    port map (
            O => \N__11282\,
            I => \N__11278\
        );

    \I__1619\ : CEMux
    port map (
            O => \N__11281\,
            I => \N__11275\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11271\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__11275\,
            I => \N__11268\
        );

    \I__1616\ : CEMux
    port map (
            O => \N__11274\,
            I => \N__11265\
        );

    \I__1615\ : Span4Mux_h
    port map (
            O => \N__11271\,
            I => \N__11262\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__11268\,
            I => \N__11259\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__11265\,
            I => \N__11256\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__11262\,
            I => \delay_measurement_inst.N_81_i_0\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__11259\,
            I => \delay_measurement_inst.N_81_i_0\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__11256\,
            I => \delay_measurement_inst.N_81_i_0\
        );

    \I__1609\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__11243\,
            I => \N__11239\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11236\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__11239\,
            I => \N__11232\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__11236\,
            I => \N__11229\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11235\,
            I => \N__11226\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__11232\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__11229\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11226\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__1599\ : InMux
    port map (
            O => \N__11219\,
            I => \bfn_5_15_0_\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__11213\,
            I => \N__11210\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__11210\,
            I => \N__11205\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11202\
        );

    \I__1594\ : InMux
    port map (
            O => \N__11208\,
            I => \N__11199\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__11205\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11202\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__11199\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__1590\ : InMux
    port map (
            O => \N__11192\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__11189\,
            I => \N__11184\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__11188\,
            I => \N__11181\
        );

    \I__1587\ : InMux
    port map (
            O => \N__11187\,
            I => \N__11178\
        );

    \I__1586\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11173\
        );

    \I__1585\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11173\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__11178\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__11173\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__1582\ : InMux
    port map (
            O => \N__11168\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__11165\,
            I => \N__11160\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__11164\,
            I => \N__11157\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11154\
        );

    \I__1578\ : InMux
    port map (
            O => \N__11160\,
            I => \N__11149\
        );

    \I__1577\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11149\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__11154\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__11149\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__1574\ : InMux
    port map (
            O => \N__11144\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__1573\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11136\
        );

    \I__1572\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11131\
        );

    \I__1571\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11131\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__11136\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__11131\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__1568\ : InMux
    port map (
            O => \N__11126\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4Z0Z_3_cascade_\
        );

    \I__1566\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__11117\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__11114\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6Z0Z_3_cascade_\
        );

    \I__1563\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__11108\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__11105\,
            I => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6_cascade_\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__11102\,
            I => \phase_controller_inst1.stoper_tr.N_92_cascade_\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__11099\,
            I => \N__11095\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__11098\,
            I => \N__11091\
        );

    \I__1557\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11087\
        );

    \I__1556\ : InMux
    port map (
            O => \N__11094\,
            I => \N__11084\
        );

    \I__1555\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11079\
        );

    \I__1554\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11079\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__11087\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__11084\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__11079\,
            I => \delay_measurement_inst.elapsed_time_tr_9\
        );

    \I__1550\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11061\
        );

    \I__1549\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11061\
        );

    \I__1548\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11049\
        );

    \I__1547\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11049\
        );

    \I__1546\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11049\
        );

    \I__1545\ : InMux
    port map (
            O => \N__11067\,
            I => \N__11049\
        );

    \I__1544\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11049\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11046\
        );

    \I__1542\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11043\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__11049\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__11046\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__11043\,
            I => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__11036\,
            I => \N__11026\
        );

    \I__1537\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11023\
        );

    \I__1536\ : InMux
    port map (
            O => \N__11034\,
            I => \N__11018\
        );

    \I__1535\ : InMux
    port map (
            O => \N__11033\,
            I => \N__11018\
        );

    \I__1534\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11007\
        );

    \I__1533\ : InMux
    port map (
            O => \N__11031\,
            I => \N__11007\
        );

    \I__1532\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11007\
        );

    \I__1531\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11007\
        );

    \I__1530\ : InMux
    port map (
            O => \N__11026\,
            I => \N__11007\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__11023\,
            I => \delay_measurement_inst.N_165\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__11018\,
            I => \delay_measurement_inst.N_165\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__11007\,
            I => \delay_measurement_inst.N_165\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__11000\,
            I => \N__10995\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__10999\,
            I => \N__10992\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__10998\,
            I => \N__10987\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10983\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10972\
        );

    \I__1521\ : InMux
    port map (
            O => \N__10991\,
            I => \N__10972\
        );

    \I__1520\ : InMux
    port map (
            O => \N__10990\,
            I => \N__10972\
        );

    \I__1519\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10972\
        );

    \I__1518\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10972\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10983\,
            I => \N__10969\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__10972\,
            I => \N__10966\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__10969\,
            I => \delay_measurement_inst.N_212\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__10966\,
            I => \delay_measurement_inst.N_212\
        );

    \I__1513\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10957\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10954\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__10957\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10954\,
            I => \delay_measurement_inst.elapsed_time_tr_4\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__10949\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10943\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__10943\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10937\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10937\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__10934\,
            I => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_15_cascade_\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10928\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__1501\ : Span12Mux_v
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1500\ : Odrv12
    port map (
            O => \N__10922\,
            I => il_max_comp2_c
        );

    \I__1499\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10916\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10916\,
            I => \il_max_comp2_D1\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10910\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__10910\,
            I => \N__10907\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__10907\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10901\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10901\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10895\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10889\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10883\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10877\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__10877\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__10871\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__10865\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10859\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10853\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\
        );

    \I__1476\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10847\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__10844\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10838\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__10829\,
            I => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__10820\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\
        );

    \I__1465\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__10811\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__10805\,
            I => \N__10802\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__10802\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10793\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10793\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\
        );

    \I__1456\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__10784\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10775\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__1450\ : InMux
    port map (
            O => \N__10772\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__10766\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10763\,
            I => \bfn_4_18_0_\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10757\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__1444\ : InMux
    port map (
            O => \N__10754\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10748\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__10748\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10745\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__10736\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10733\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10730\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__1435\ : CEMux
    port map (
            O => \N__10727\,
            I => \N__10712\
        );

    \I__1434\ : CEMux
    port map (
            O => \N__10726\,
            I => \N__10712\
        );

    \I__1433\ : CEMux
    port map (
            O => \N__10725\,
            I => \N__10712\
        );

    \I__1432\ : CEMux
    port map (
            O => \N__10724\,
            I => \N__10712\
        );

    \I__1431\ : CEMux
    port map (
            O => \N__10723\,
            I => \N__10712\
        );

    \I__1430\ : GlobalMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__1429\ : gio2CtrlBuf
    port map (
            O => \N__10709\,
            I => \delay_measurement_inst.delay_tr_timer.N_138_i_g\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__10703\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__10697\,
            I => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10694\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10691\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10688\,
            I => \bfn_4_17_0_\
        );

    \I__1421\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__10682\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10679\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__1418\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10673\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10670\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__1415\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10664\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10661\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__1412\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10655\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__10655\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10652\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10646\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10643\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__1406\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__10637\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__1404\ : InMux
    port map (
            O => \N__10634\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10631\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10621\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__1399\ : Odrv12
    port map (
            O => \N__10621\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__10618\,
            I => \delay_measurement_inst.elapsed_time_tr_10\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10613\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10606\
        );

    \I__1395\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10603\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10606\,
            I => \N__10600\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__10603\,
            I => \N__10597\
        );

    \I__1392\ : Odrv12
    port map (
            O => \N__10600\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__10597\,
            I => \delay_measurement_inst.elapsed_time_tr_11\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10592\,
            I => \bfn_4_16_0_\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10585\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10582\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10585\,
            I => \N__10579\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__10582\,
            I => \N__10576\
        );

    \I__1385\ : Odrv12
    port map (
            O => \N__10579\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__10576\,
            I => \delay_measurement_inst.elapsed_time_tr_12\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10571\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__1382\ : InMux
    port map (
            O => \N__10568\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10556\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10556\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10553\
        );

    \I__1378\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10550\
        );

    \I__1377\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10547\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__10556\,
            I => \N__10544\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10553\,
            I => \N__10537\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10550\,
            I => \N__10537\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__10547\,
            I => \N__10537\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__10544\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__10537\,
            I => \delay_measurement_inst.elapsed_time_tr_14\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10532\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__10529\,
            I => \N__10525\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__10528\,
            I => \N__10521\
        );

    \I__1367\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10513\
        );

    \I__1366\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10513\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10510\
        );

    \I__1364\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10505\
        );

    \I__1363\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10505\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10502\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__10513\,
            I => \N__10499\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10492\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10492\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__10502\,
            I => \N__10492\
        );

    \I__1357\ : Span4Mux_h
    port map (
            O => \N__10499\,
            I => \N__10489\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__10492\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__10489\,
            I => \delay_measurement_inst.elapsed_time_tr_15\
        );

    \I__1354\ : InMux
    port map (
            O => \N__10484\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10473\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10468\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10468\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10463\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__10468\,
            I => \N__10463\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__10463\,
            I => \delay_measurement_inst.elapsed_time_tr_16\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10460\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__10457\,
            I => \N__10452\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__10456\,
            I => \N__10449\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10443\
        );

    \I__1342\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10443\
        );

    \I__1341\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10440\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10437\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10443\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__10440\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__10437\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\
        );

    \I__1336\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__10427\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_3\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10420\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10417\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10420\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10417\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10408\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10405\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10401\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10398\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10395\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__10401\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__10398\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10395\,
            I => \delay_measurement_inst.elapsed_time_tr_3\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10388\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__1321\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10378\
        );

    \I__1319\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10375\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__10378\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__10375\,
            I => \delay_measurement_inst.elapsed_time_tr_5\
        );

    \I__1316\ : InMux
    port map (
            O => \N__10370\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10357\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__10360\,
            I => \N__10354\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__10357\,
            I => \N__10350\
        );

    \I__1310\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10347\
        );

    \I__1309\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10344\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__10350\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__10347\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10344\,
            I => \delay_measurement_inst.elapsed_time_tr_6\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10337\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10331\,
            I => \N__10326\
        );

    \I__1302\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10323\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10320\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__10326\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__10323\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10320\,
            I => \delay_measurement_inst.elapsed_time_tr_7\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10313\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__10304\,
            I => \N__10299\
        );

    \I__1293\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10296\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10293\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__10299\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__10296\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__10293\,
            I => \delay_measurement_inst.elapsed_time_tr_8\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10286\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__10283\,
            I => \N__10279\
        );

    \I__1286\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10274\
        );

    \I__1285\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10274\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__10274\,
            I => \delay_measurement_inst.N_200\
        );

    \I__1283\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__10268\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_3\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__10265\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\
        );

    \I__1280\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10259\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__10259\,
            I => \delay_measurement_inst.un1_tr_state_1_i_0_a2_0_7\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10250\
        );

    \I__1277\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10250\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__10250\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__10247\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10241\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__10241\,
            I => \delay_measurement_inst.delay_tr_timer.N_203\
        );

    \I__1272\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__10235\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\
        );

    \I__1270\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10228\
        );

    \I__1269\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10222\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__10225\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__10222\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__1265\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__10214\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\
        );

    \I__1263\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10207\
        );

    \I__1262\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10204\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__10207\,
            I => \N__10201\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__10204\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__10201\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10193\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__10193\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\
        );

    \I__1256\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10186\
        );

    \I__1255\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10186\,
            I => \N__10180\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__10183\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__10180\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__1251\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__10172\,
            I => \delay_measurement_inst.N_168\
        );

    \I__1249\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10163\
        );

    \I__1248\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10163\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__10163\,
            I => \delay_measurement_inst.N_81_i\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__10160\,
            I => \delay_measurement_inst.N_81_i_cascade_\
        );

    \I__1245\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10153\
        );

    \I__1244\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10149\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__10153\,
            I => \N__10146\
        );

    \I__1242\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10143\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__10149\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__10146\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__10143\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__1238\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__10133\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__10130\,
            I => \N__10127\
        );

    \I__1235\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10124\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__10124\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\
        );

    \I__1233\ : InMux
    port map (
            O => \N__10121\,
            I => \N__10118\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10118\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\
        );

    \I__1231\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10111\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10108\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__10111\,
            I => \N__10105\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__10108\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__10105\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__1226\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10097\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__10097\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\
        );

    \I__1224\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10090\
        );

    \I__1223\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10087\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10090\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__10087\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__1220\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__10079\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\
        );

    \I__1218\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10072\
        );

    \I__1217\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10066\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__10069\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__10066\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__1213\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10058\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10058\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\
        );

    \I__1211\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10051\
        );

    \I__1210\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10048\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__10051\,
            I => \N__10045\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__10048\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__10045\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__1206\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__10037\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\
        );

    \I__1204\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10030\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10027\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__10030\,
            I => \N__10024\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__10027\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__10024\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__1199\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__10016\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\
        );

    \I__1197\ : InMux
    port map (
            O => \N__10013\,
            I => \N__10009\
        );

    \I__1196\ : InMux
    port map (
            O => \N__10012\,
            I => \N__10006\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__10009\,
            I => \N__10003\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__10006\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__10003\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9992\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9992\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_13\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9983\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_14\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__9974\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_15\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9965\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__9965\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_16\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__9962\,
            I => \N__9959\
        );

    \I__1179\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9956\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_17\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1176\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9947\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__9947\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_18\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9938\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__9938\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_19\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9935\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__9932\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__1168\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9923\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__9923\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\
        );

    \I__1166\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9917\,
            I => \N__9913\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9910\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__9913\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__9910\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1160\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__9899\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_5\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9892\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9889\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9892\,
            I => \N__9886\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9889\,
            I => \N__9883\
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__9886\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__9883\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9872\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_6\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9866\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__9866\,
            I => \N__9862\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9859\
        );

    \I__1146\ : Odrv12
    port map (
            O => \N__9862\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9859\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__9854\,
            I => \N__9851\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9848\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_7\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__9845\,
            I => \N__9842\
        );

    \I__1140\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9838\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9841\,
            I => \N__9835\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__9838\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9835\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__9830\,
            I => \N__9827\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9824\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_8\
        );

    \I__1133\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9814\
        );

    \I__1131\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9811\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__9814\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9811\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__9806\,
            I => \N__9803\
        );

    \I__1127\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9800\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__9800\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_9\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9794\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9794\,
            I => \N__9790\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__9790\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__9787\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__9782\,
            I => \N__9779\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9776\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9776\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_10\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9767\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9767\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_11\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__9764\,
            I => \N__9761\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9758\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_12\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__9755\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19_cascade_\
        );

    \I__1110\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__9749\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9743\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__9743\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__9740\,
            I => \N__9737\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9734\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9734\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_1\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__9728\,
            I => \N__9724\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9721\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__9724\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__9721\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__9716\,
            I => \N__9713\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__9710\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_2\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__9704\,
            I => \N__9700\
        );

    \I__1093\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9697\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__9700\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9697\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9686\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9686\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_3\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9680\,
            I => \N__9676\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__1084\ : Odrv12
    port map (
            O => \N__9676\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__9673\,
            I => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__9662\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_i_4\
        );

    \I__1079\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9656\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__9656\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__9650\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9644\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__9644\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9638\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__9638\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9632\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__9629\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9623\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__9623\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__9617\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\
        );

    \I__1064\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9611\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9611\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__9608\,
            I => \N__9605\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9601\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9598\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__9601\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__9598\,
            I => \delay_measurement_inst.elapsed_time_tr_1\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9586\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9586\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9583\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9586\,
            I => \N__9580\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9583\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__9580\,
            I => \delay_measurement_inst.elapsed_time_tr_2\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9572\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__9569\,
            I => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5_cascade_\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9563\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9557\,
            I => \N__9554\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__9554\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__9545\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9539\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9533\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9530\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__9530\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__9527\,
            I => \delay_measurement_inst.N_212_cascade_\
        );

    \I__1034\ : InMux
    port map (
            O => \N__9524\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9521\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9518\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9515\,
            I => \bfn_2_24_0_\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9512\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9509\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9503\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__9500\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9497\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__9488\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9485\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9479\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__9479\,
            I => \N__9476\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__9476\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9473\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__9470\,
            I => \N__9467\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__9464\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9461\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__9452\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\
        );

    \I__1009\ : InMux
    port map (
            O => \N__9449\,
            I => \bfn_2_23_0_\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__9437\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9434\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9431\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9428\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9425\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__9416\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\
        );

    \I__997\ : InMux
    port map (
            O => \N__9413\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\
        );

    \I__996\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__9404\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\
        );

    \I__993\ : InMux
    port map (
            O => \N__9401\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\
        );

    \I__992\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__990\ : Odrv4
    port map (
            O => \N__9392\,
            I => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\
        );

    \I__989\ : InMux
    port map (
            O => \N__9389\,
            I => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\
        );

    \I__988\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9383\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__9383\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\
        );

    \I__986\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9376\
        );

    \I__985\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9373\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9370\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9373\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__982\ : Odrv4
    port map (
            O => \N__9370\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__980\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9359\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\
        );

    \I__978\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9352\
        );

    \I__977\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9349\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__9352\,
            I => \N__9346\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__9349\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__9346\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__973\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9338\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\
        );

    \I__971\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9331\
        );

    \I__970\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9325\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__9328\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__9325\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__966\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9317\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\
        );

    \I__964\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9310\
        );

    \I__963\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__9307\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__9304\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__9299\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\
        );

    \I__958\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9293\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\
        );

    \I__956\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__9287\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\
        );

    \I__954\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9280\
        );

    \I__953\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9277\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9280\,
            I => \N__9274\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9277\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__9274\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__949\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__9266\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\
        );

    \I__947\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9259\
        );

    \I__946\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9256\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9259\,
            I => \N__9253\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9256\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__9253\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__941\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__9242\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\
        );

    \I__939\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9235\
        );

    \I__938\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9232\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__9232\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__9229\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__934\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__9221\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\
        );

    \I__932\ : InMux
    port map (
            O => \N__9218\,
            I => \N__9214\
        );

    \I__931\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9208\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__9211\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__9208\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__926\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__9197\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\
        );

    \I__924\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9190\
        );

    \I__923\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9187\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__9187\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__9184\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__919\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9176\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\
        );

    \I__917\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9169\
        );

    \I__916\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9169\,
            I => \N__9163\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__9166\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__913\ : Odrv4
    port map (
            O => \N__9163\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__911\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__9152\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\
        );

    \I__909\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9145\
        );

    \I__908\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9142\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__9142\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__905\ : Odrv4
    port map (
            O => \N__9139\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__903\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__9128\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_13\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9122\
        );

    \I__900\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__9119\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_14\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__897\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__9110\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_15\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__894\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__9101\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_16\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__891\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9092\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__9092\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_17\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__888\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__9083\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_18\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__885\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__9074\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_19\
        );

    \I__883\ : InMux
    port map (
            O => \N__9071\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__882\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__9065\,
            I => \N__9062\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__9062\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\
        );

    \I__879\ : InMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__9056\,
            I => \N__9052\
        );

    \I__877\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9049\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__9052\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__9049\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__873\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__9038\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_5\
        );

    \I__871\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__9032\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\
        );

    \I__869\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__9022\
        );

    \I__867\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9019\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__9022\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__9019\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__863\ : InMux
    port map (
            O => \N__9011\,
            I => \N__9008\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__9008\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_6\
        );

    \I__861\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8998\
        );

    \I__859\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8995\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__8998\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8995\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__8990\,
            I => \N__8987\
        );

    \I__855\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8984\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__8984\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_7\
        );

    \I__853\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8974\
        );

    \I__851\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8971\
        );

    \I__850\ : Odrv12
    port map (
            O => \N__8974\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__8971\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__8966\,
            I => \N__8963\
        );

    \I__847\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8960\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_8\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__8957\,
            I => \N__8954\
        );

    \I__844\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8951\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__8951\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_9\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__841\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__8942\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_10\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__838\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__8933\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_11\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__8930\,
            I => \N__8927\
        );

    \I__835\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__8924\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_12\
        );

    \I__833\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8918\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__830\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8908\
        );

    \I__829\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8904\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8901\
        );

    \I__827\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8898\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8904\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__8901\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8898\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__822\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__8885\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_1\
        );

    \I__820\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8879\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8879\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\
        );

    \I__818\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8869\
        );

    \I__816\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__8869\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__8866\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__812\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8855\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_2\
        );

    \I__810\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__8849\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\
        );

    \I__808\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8843\,
            I => \N__8839\
        );

    \I__806\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8836\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__8839\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8836\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__802\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8825\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_3\
        );

    \I__800\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__8816\,
            I => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\
        );

    \I__797\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8810\,
            I => \N__8806\
        );

    \I__795\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8803\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__8806\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8803\,
            I => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__791\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8792\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_i_4\
        );

    \I__789\ : InMux
    port map (
            O => \N__8789\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\
        );

    \I__788\ : InMux
    port map (
            O => \N__8786\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\
        );

    \I__787\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__8780\,
            I => \N_27_i_i\
        );

    \I__785\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8774\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8774\,
            I => un7_start_stop
        );

    \I__783\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__8768\,
            I => \N__8765\
        );

    \I__781\ : Span12Mux_s5_v
    port map (
            O => \N__8765\,
            I => \N__8762\
        );

    \I__780\ : Span12Mux_h
    port map (
            O => \N__8762\,
            I => \N__8759\
        );

    \I__779\ : Span12Mux_h
    port map (
            O => \N__8759\,
            I => \N__8753\
        );

    \I__778\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8750\
        );

    \I__777\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8747\
        );

    \I__776\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8744\
        );

    \I__775\ : Odrv12
    port map (
            O => \N__8753\,
            I => \CONSTANT_ONE_NET\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8750\,
            I => \CONSTANT_ONE_NET\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__8747\,
            I => \CONSTANT_ONE_NET\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8744\,
            I => \CONSTANT_ONE_NET\
        );

    \I__771\ : InMux
    port map (
            O => \N__8735\,
            I => \bfn_1_19_0_\
        );

    \I__770\ : InMux
    port map (
            O => \N__8732\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\
        );

    \I__769\ : InMux
    port map (
            O => \N__8729\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\
        );

    \I__768\ : InMux
    port map (
            O => \N__8726\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\
        );

    \I__767\ : InMux
    port map (
            O => \N__8723\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\
        );

    \I__766\ : InMux
    port map (
            O => \N__8720\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\
        );

    \I__765\ : InMux
    port map (
            O => \N__8717\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\
        );

    \I__764\ : InMux
    port map (
            O => \N__8714\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\
        );

    \I__763\ : InMux
    port map (
            O => \N__8711\,
            I => \bfn_1_20_0_\
        );

    \I__762\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__8702\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\
        );

    \I__759\ : InMux
    port map (
            O => \N__8699\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__757\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__8690\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\
        );

    \I__755\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__8681\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\
        );

    \I__752\ : InMux
    port map (
            O => \N__8678\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\
        );

    \I__751\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__8669\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\
        );

    \I__748\ : InMux
    port map (
            O => \N__8666\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\
        );

    \I__747\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__8657\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\
        );

    \I__744\ : InMux
    port map (
            O => \N__8654\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\
        );

    \I__743\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__8645\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\
        );

    \I__740\ : InMux
    port map (
            O => \N__8642\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\
        );

    \I__739\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8636\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__737\ : Odrv4
    port map (
            O => \N__8633\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\
        );

    \I__736\ : InMux
    port map (
            O => \N__8630\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\
        );

    \I__735\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__8621\,
            I => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\
        );

    \I__732\ : InMux
    port map (
            O => \N__8618\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\
        );

    \I__731\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8612\,
            I => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0\
        );

    \IN_MUX_bfv_1_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_18_0_\
        );

    \IN_MUX_bfv_1_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_1_19_0_\
        );

    \IN_MUX_bfv_1_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_1_20_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_3_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_3_21_0_\
        );

    \IN_MUX_bfv_2_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_22_0_\
        );

    \IN_MUX_bfv_2_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_2_23_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_7_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_7_21_0_\
        );

    \IN_MUX_bfv_9_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_17_0_\
        );

    \IN_MUX_bfv_9_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            carryinitout => \bfn_9_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_2_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_2_17_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_4_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_4_17_0_\
        );

    \IN_MUX_bfv_4_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_4_18_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_5_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_5_17_0_\
        );

    \IN_MUX_bfv_5_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_5_18_0_\
        );

    \IN_MUX_bfv_8_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_26_0_\
        );

    \IN_MUX_bfv_8_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_27_0_\
        );

    \IN_MUX_bfv_8_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_28_0_\
        );

    \IN_MUX_bfv_8_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_29_0_\
        );

    \IN_MUX_bfv_9_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_26_0_\
        );

    \IN_MUX_bfv_9_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_9_27_0_\
        );

    \IN_MUX_bfv_9_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_9_28_0_\
        );

    \IN_MUX_bfv_9_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_9_29_0_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19511\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_138_i_g\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21734\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_hc_timer.N_136_i_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__8756\,
            CLKHFEN => \N__8758\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__8757\,
            RGB2PWM => \N__8783\,
            RGB1 => rgb_g_wire,
            CURREN => \N__8771\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__8777\,
            RGB0PWM => \N__22342\,
            RGB0 => rgb_r_wire
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__21458\,
            GLOBALBUFFEROUTPUT => \delay_measurement_inst.delay_tr_timer.N_139_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_0_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15111\,
            in1 => \N__15069\,
            in2 => \N__19907\,
            in3 => \N__15170\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22041\,
            ce => \N__21315\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_8_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15064\,
            in1 => \N__19860\,
            in2 => \N__15262\,
            in3 => \N__8627\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_1_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15254\,
            in1 => \N__15065\,
            in2 => \N__19898\,
            in3 => \N__8615\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_5_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15062\,
            in1 => \N__19858\,
            in2 => \N__15260\,
            in3 => \N__8663\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_7_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15257\,
            in1 => \N__15068\,
            in2 => \N__19901\,
            in3 => \N__8639\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_3_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15061\,
            in1 => \N__19857\,
            in2 => \N__15259\,
            in3 => \N__8687\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_2_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15255\,
            in1 => \N__15066\,
            in2 => \N__19899\,
            in3 => \N__8708\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_6_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15063\,
            in1 => \N__19859\,
            in2 => \N__15261\,
            in3 => \N__8651\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_4_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15256\,
            in1 => \N__15067\,
            in2 => \N__19900\,
            in3 => \N__8675\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22036\,
            ce => 'H',
            sr => \N__22278\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_1_LC_1_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__15102\,
            in1 => \_gnd_net_\,
            in2 => \N__14953\,
            in3 => \N__8911\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1B6_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14946\,
            in2 => \_gnd_net_\,
            in3 => \N__15101\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_RNIG1BZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_1_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9296\,
            in2 => \N__8915\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_18_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8876\,
            in2 => \_gnd_net_\,
            in3 => \N__8699\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_3_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8846\,
            in2 => \N__8696\,
            in3 => \N__8678\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_4_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8813\,
            in2 => \_gnd_net_\,
            in3 => \N__8666\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_5_LC_1_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9059\,
            in2 => \_gnd_net_\,
            in3 => \N__8654\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_6_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9029\,
            in2 => \_gnd_net_\,
            in3 => \N__8642\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_7_LC_1_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9005\,
            in2 => \_gnd_net_\,
            in3 => \N__8630\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_8_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8981\,
            in2 => \_gnd_net_\,
            in3 => \N__8618\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_9_LC_1_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9148\,
            in2 => \_gnd_net_\,
            in3 => \N__8735\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_9\,
            ltout => OPEN,
            carryin => \bfn_1_19_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_10_LC_1_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9193\,
            in2 => \_gnd_net_\,
            in3 => \N__8732\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_11_LC_1_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9172\,
            in2 => \_gnd_net_\,
            in3 => \N__8729\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_12_LC_1_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9262\,
            in2 => \_gnd_net_\,
            in3 => \N__8726\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_13_LC_1_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9217\,
            in2 => \_gnd_net_\,
            in3 => \N__8723\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_14_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9379\,
            in2 => \_gnd_net_\,
            in3 => \N__8720\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_15_LC_1_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9283\,
            in2 => \_gnd_net_\,
            in3 => \N__8717\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_16_LC_1_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9238\,
            in2 => \_gnd_net_\,
            in3 => \N__8714\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_17_LC_1_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9313\,
            in2 => \_gnd_net_\,
            in3 => \N__8711\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_17\,
            ltout => OPEN,
            carryin => \bfn_1_20_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_18_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9355\,
            in2 => \_gnd_net_\,
            in3 => \N__8789\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_19_LC_1_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9334\,
            in2 => \_gnd_net_\,
            in3 => \N__8786\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_RNO_0_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \reset_ibuf_gb_io_RNI79U7_LC_1_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => red_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.N_27_i_i_LC_1_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21721\,
            in2 => \_gnd_net_\,
            in3 => \N__22340\,
            lcout => \N_27_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un7_start_stop_LC_1_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22341\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21725\,
            lcout => un7_start_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11249\,
            lcout => \delay_measurement_inst.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22042\,
            ce => \N__10727\,
            sr => \N__22254\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11216\,
            lcout => \delay_measurement_inst.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22042\,
            ce => \N__10727\,
            sr => \N__22254\
        );

    \phase_controller_slave.stoper_tr.target_time_2_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__13266\,
            in1 => \N__13327\,
            in2 => \N__13307\,
            in3 => \N__13354\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22038\,
            ce => \N__13823\,
            sr => \N__22260\
        );

    \phase_controller_slave.stoper_tr.target_time_4_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__20135\,
            in1 => \N__13231\,
            in2 => \N__12857\,
            in3 => \N__13155\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22038\,
            ce => \N__13823\,
            sr => \N__22260\
        );

    \phase_controller_slave.stoper_tr.target_time_5_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__13156\,
            in1 => \N__12738\,
            in2 => \N__13235\,
            in3 => \N__20136\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22038\,
            ce => \N__13823\,
            sr => \N__22260\
        );

    \phase_controller_slave.stoper_tr.target_time_1_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__12712\,
            in1 => \N__13302\,
            in2 => \N__12700\,
            in3 => \N__13267\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22038\,
            ce => \N__13823\,
            sr => \N__22260\
        );

    \phase_controller_slave.stoper_tr.target_time_3_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__13326\,
            in1 => \N__13306\,
            in2 => \_gnd_net_\,
            in3 => \N__13268\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22038\,
            ce => \N__13823\,
            sr => \N__22260\
        );

    \phase_controller_slave.stoper_tr.target_time_6_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110001"
        )
    port map (
            in0 => \N__13157\,
            in1 => \N__20137\,
            in2 => \N__13183\,
            in3 => \N__13232\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22038\,
            ce => \N__13823\,
            sr => \N__22260\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8921\,
            in2 => \N__8891\,
            in3 => \N__8907\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8882\,
            in2 => \N__8861\,
            in3 => \N__8872\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8852\,
            in2 => \N__8831\,
            in3 => \N__8842\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8822\,
            in2 => \N__8798\,
            in3 => \N__8809\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9068\,
            in2 => \N__9044\,
            in3 => \N__9055\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9035\,
            in2 => \N__9014\,
            in3 => \N__9025\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9659\,
            in2 => \N__8990\,
            in3 => \N__9001\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9536\,
            in2 => \N__8966\,
            in3 => \N__8977\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9566\,
            in2 => \N__8957\,
            in3 => \N__9149\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_2_16_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9542\,
            in2 => \N__8948\,
            in3 => \N__9194\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9653\,
            in2 => \N__8939\,
            in3 => \N__9173\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9560\,
            in2 => \N__8930\,
            in3 => \N__9263\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9551\,
            in2 => \N__9134\,
            in3 => \N__9218\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9614\,
            in2 => \N__9125\,
            in3 => \N__9380\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9626\,
            in2 => \N__9116\,
            in3 => \N__9284\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9635\,
            in2 => \N__9107\,
            in3 => \N__9239\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_2_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9620\,
            in2 => \N__9098\,
            in3 => \N__9314\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_2_17_0_\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_2_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9641\,
            in2 => \N__9089\,
            in3 => \N__9356\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9647\,
            in2 => \N__9080\,
            in3 => \N__9335\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_2_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9071\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_slave.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9299\,
            in3 => \N__14945\,
            lcout => \phase_controller_slave.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNI38A6_0_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__15171\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15002\,
            lcout => \phase_controller_slave.stoper_tr.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_15_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__15071\,
            in1 => \N__19892\,
            in2 => \N__15263\,
            in3 => \N__9290\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_12_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15228\,
            in1 => \N__15075\,
            in2 => \N__19904\,
            in3 => \N__9269\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_16_LC_2_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15072\,
            in1 => \N__19893\,
            in2 => \N__9248\,
            in3 => \N__15232\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_13_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15229\,
            in1 => \N__15076\,
            in2 => \N__19905\,
            in3 => \N__9224\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_10_LC_2_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15070\,
            in1 => \N__19891\,
            in2 => \N__9203\,
            in3 => \N__15231\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_11_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15227\,
            in1 => \N__15074\,
            in2 => \N__19903\,
            in3 => \N__9179\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_9_LC_2_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__15073\,
            in1 => \N__19894\,
            in2 => \N__9158\,
            in3 => \N__15233\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_14_LC_2_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15230\,
            in1 => \N__15077\,
            in2 => \N__19906\,
            in3 => \N__9386\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22026\,
            ce => 'H',
            sr => \N__22284\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_18_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__15235\,
            in1 => \N__19878\,
            in2 => \N__9365\,
            in3 => \N__15079\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22022\,
            ce => 'H',
            sr => \N__22289\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_19_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__15078\,
            in1 => \N__15236\,
            in2 => \N__19902\,
            in3 => \N__9341\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22022\,
            ce => 'H',
            sr => \N__22289\
        );

    \phase_controller_slave.stoper_tr.accumulated_time_17_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__15234\,
            in1 => \N__19877\,
            in2 => \N__15083\,
            in3 => \N__9320\,
            lcout => \phase_controller_slave.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22022\,
            ce => 'H',
            sr => \N__22289\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_4_LC_2_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12354\,
            in1 => \N__15651\,
            in2 => \N__12499\,
            in3 => \N__9398\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_6_LC_2_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12484\,
            in1 => \N__12358\,
            in2 => \N__15701\,
            in3 => \N__9494\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_2_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12353\,
            in1 => \N__15650\,
            in2 => \N__12498\,
            in3 => \N__9422\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_1_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12482\,
            in1 => \N__12356\,
            in2 => \N__15699\,
            in3 => \N__10136\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_5_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12355\,
            in1 => \N__15652\,
            in2 => \N__12500\,
            in3 => \N__9506\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_3_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12483\,
            in1 => \N__12357\,
            in2 => \N__15700\,
            in3 => \N__9410\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_7_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12485\,
            in1 => \N__12359\,
            in2 => \N__15702\,
            in3 => \N__9482\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22018\,
            ce => 'H',
            sr => \N__22293\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_10_LC_2_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__12479\,
            in1 => \N__15729\,
            in2 => \N__9446\,
            in3 => \N__12351\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22013\,
            ce => 'H',
            sr => \N__22297\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_9_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12350\,
            in1 => \N__12481\,
            in2 => \N__15737\,
            in3 => \N__9458\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22013\,
            ce => 'H',
            sr => \N__22297\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_8_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__12480\,
            in1 => \N__15730\,
            in2 => \N__9470\,
            in3 => \N__12352\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22013\,
            ce => 'H',
            sr => \N__22297\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10157\,
            in2 => \N__9929\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_22_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_2_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9731\,
            in2 => \_gnd_net_\,
            in3 => \N__9413\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_3_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9707\,
            in2 => \N__10130\,
            in3 => \N__9401\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_4_LC_2_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9683\,
            in2 => \_gnd_net_\,
            in3 => \N__9389\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_5_LC_2_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9920\,
            in2 => \_gnd_net_\,
            in3 => \N__9497\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_6_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9896\,
            in2 => \_gnd_net_\,
            in3 => \N__9485\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_7_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9869\,
            in2 => \_gnd_net_\,
            in3 => \N__9473\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_8_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9845\,
            in3 => \N__9461\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_8\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_9_LC_2_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9821\,
            in2 => \_gnd_net_\,
            in3 => \N__9449\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_9\,
            ltout => OPEN,
            carryin => \bfn_2_23_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_10_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9797\,
            in2 => \_gnd_net_\,
            in3 => \N__9434\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_11_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10114\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_12_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10012\,
            in2 => \_gnd_net_\,
            in3 => \N__9428\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_13_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10075\,
            in2 => \_gnd_net_\,
            in3 => \N__9425\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_14_LC_2_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10033\,
            in2 => \_gnd_net_\,
            in3 => \N__9524\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_15_LC_2_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10054\,
            in2 => \_gnd_net_\,
            in3 => \N__9521\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_16_LC_2_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10094\,
            in2 => \_gnd_net_\,
            in3 => \N__9518\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_16\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_17_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10210\,
            in2 => \_gnd_net_\,
            in3 => \N__9515\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_17\,
            ltout => OPEN,
            carryin => \bfn_2_24_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_18_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10189\,
            in2 => \_gnd_net_\,
            in3 => \N__9512\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_19_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10231\,
            in2 => \_gnd_net_\,
            in3 => \N__9509\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_8_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__11034\,
            in1 => \N__10169\,
            in2 => \N__12776\,
            in3 => \N__10310\,
            lcout => measured_delay_tr_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22043\,
            ce => 'H',
            sr => \N__22242\
        );

    \delay_measurement_inst.delay_tr_reg_7_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__11033\,
            in1 => \N__10168\,
            in2 => \N__12817\,
            in3 => \N__10334\,
            lcout => measured_delay_tr_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22043\,
            ce => 'H',
            sr => \N__22242\
        );

    \delay_measurement_inst.delay_tr_reg_esr_5_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__11067\,
            in1 => \N__11029\,
            in2 => \N__10998\,
            in3 => \N__10385\,
            lcout => measured_delay_tr_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_esr_2_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__9591\,
            in1 => \N__10986\,
            in2 => \N__11036\,
            in3 => \N__11066\,
            lcout => measured_delay_tr_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_esr_16_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__11364\,
            in1 => \_gnd_net_\,
            in2 => \N__10481\,
            in3 => \N__20940\,
            lcout => measured_delay_tr_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_ess_1_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__11031\,
            in1 => \N__10991\,
            in2 => \N__9608\,
            in3 => \N__11069\,
            lcout => measured_delay_tr_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_esr_15_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__11363\,
            in1 => \N__10282\,
            in2 => \N__10528\,
            in3 => \N__20942\,
            lcout => measured_delay_tr_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_esr_14_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__20941\,
            in1 => \N__10563\,
            in2 => \N__10283\,
            in3 => \N__11362\,
            lcout => measured_delay_tr_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_ess_3_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__11070\,
            in1 => \N__11032\,
            in2 => \N__10999\,
            in3 => \N__10412\,
            lcout => measured_delay_tr_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \delay_measurement_inst.delay_tr_reg_esr_6_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__10990\,
            in2 => \N__10367\,
            in3 => \N__11068\,
            lcout => measured_delay_tr_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22039\,
            ce => \N__11274\,
            sr => \N__22248\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_13_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__20070\,
            in1 => \N__19996\,
            in2 => \_gnd_net_\,
            in3 => \N__12952\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI43GB_6_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10302\,
            in1 => \N__10329\,
            in2 => \_gnd_net_\,
            in3 => \N__10353\,
            lcout => \delay_measurement_inst.N_212\,
            ltout => \delay_measurement_inst.N_212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIC9OF1_14_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10524\,
            in1 => \N__10561\,
            in2 => \N__9527\,
            in3 => \N__10423\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2_1_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13325\,
            in2 => \_gnd_net_\,
            in3 => \N__13353\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_o2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4T357_15_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__11361\,
            in1 => \_gnd_net_\,
            in2 => \N__10529\,
            in3 => \N__10256\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNI4T357_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6FAF_1_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9592\,
            in1 => \N__9604\,
            in2 => \N__10360\,
            in3 => \N__11090\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ5M42_2_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__10404\,
            in1 => \N__9593\,
            in2 => \N__11098\,
            in3 => \N__10430\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_2_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10255\,
            in1 => \N__9575\,
            in2 => \N__9569\,
            in3 => \N__11360\,
            lcout => \delay_measurement_inst.N_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.target_time_9_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011110101"
        )
    port map (
            in0 => \N__12906\,
            in1 => \N__20020\,
            in2 => \N__12586\,
            in3 => \N__12544\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_12_LC_3_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13019\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_13_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12905\,
            in2 => \_gnd_net_\,
            in3 => \N__12994\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_10_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__12881\,
            in1 => \_gnd_net_\,
            in2 => \N__12910\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_8_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__13154\,
            in1 => \_gnd_net_\,
            in2 => \N__20131\,
            in3 => \N__12777\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_7_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12818\,
            in1 => \N__20109\,
            in2 => \_gnd_net_\,
            in3 => \N__13153\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_11_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12903\,
            in2 => \_gnd_net_\,
            in3 => \N__12611\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22035\,
            ce => \N__13822\,
            sr => \N__22261\
        );

    \phase_controller_slave.stoper_tr.target_time_19_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13783\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22031\,
            ce => \N__13812\,
            sr => \N__22270\
        );

    \phase_controller_slave.stoper_tr.target_time_18_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13690\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22031\,
            ce => \N__13812\,
            sr => \N__22270\
        );

    \phase_controller_slave.stoper_tr.target_time_16_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13648\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22031\,
            ce => \N__13812\,
            sr => \N__22270\
        );

    \phase_controller_slave.stoper_tr.target_time_15_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20130\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22031\,
            ce => \N__13812\,
            sr => \N__22270\
        );

    \phase_controller_slave.stoper_tr.target_time_17_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13732\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22031\,
            ce => \N__13812\,
            sr => \N__22270\
        );

    \phase_controller_slave.stoper_tr.target_time_14_LC_3_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__20019\,
            in1 => \N__20129\,
            in2 => \_gnd_net_\,
            in3 => \N__12961\,
            lcout => \phase_controller_slave.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22031\,
            ce => \N__13812\,
            sr => \N__22270\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10640\,
            in1 => \N__10649\,
            in2 => \N__10781\,
            in3 => \N__10658\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_6_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10667\,
            in2 => \_gnd_net_\,
            in3 => \N__10676\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_0_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10685\,
            in1 => \N__9746\,
            in2 => \N__9755\,
            in3 => \N__9752\,
            lcout => \delay_measurement_inst.elapsed_time_ns_1_RNIBSKT4_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10751\,
            in1 => \N__10760\,
            in2 => \N__10742\,
            in3 => \N__10769\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr_reg_7_i_o2_7_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0_c_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10841\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10850\,
            in2 => \N__9740\,
            in3 => \N__10152\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10856\,
            in2 => \N__9716\,
            in3 => \N__9727\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10700\,
            in2 => \N__9692\,
            in3 => \N__9703\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10826\,
            in2 => \N__9668\,
            in3 => \N__9679\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10706\,
            in2 => \N__9905\,
            in3 => \N__9916\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10835\,
            in2 => \N__9878\,
            in3 => \N__9895\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10862\,
            in2 => \N__9854\,
            in3 => \N__9865\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10913\,
            in2 => \N__9830\,
            in3 => \N__9841\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10892\,
            in2 => \N__9806\,
            in3 => \N__9817\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10808\,
            in2 => \N__9782\,
            in3 => \N__9793\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10790\,
            in2 => \N__9773\,
            in3 => \N__10115\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10817\,
            in2 => \N__9764\,
            in3 => \N__10013\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10799\,
            in2 => \N__9998\,
            in3 => \N__10076\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10898\,
            in2 => \N__9989\,
            in3 => \N__10034\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10904\,
            in2 => \N__9980\,
            in3 => \N__10055\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_3_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10093\,
            in1 => \N__10874\,
            in2 => \N__9971\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_3_21_0_\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_3_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10868\,
            in2 => \N__9962\,
            in3 => \N__10211\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_3_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10880\,
            in2 => \N__9953\,
            in3 => \N__10190\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_3_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10886\,
            in2 => \N__9944\,
            in3 => \N__10232\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_3_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9935\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9932\,
            in3 => \N__18101\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_RNO_0_1_LC_3_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__18051\,
            in1 => \_gnd_net_\,
            in2 => \N__18109\,
            in3 => \N__10156\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSR_LC_3_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18102\,
            in2 => \_gnd_net_\,
            in3 => \N__18050\,
            lcout => \phase_controller_slave.stoper_hc.un1_accumulated_time_cry_19_c_RNIVGSRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_11_LC_3_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12467\,
            in1 => \N__12347\,
            in2 => \N__15734\,
            in3 => \N__10121\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22000\,
            ce => 'H',
            sr => \N__22298\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_16_LC_3_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12346\,
            in1 => \N__15716\,
            in2 => \N__12497\,
            in3 => \N__10100\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22000\,
            ce => 'H',
            sr => \N__22298\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_13_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12468\,
            in1 => \N__12348\,
            in2 => \N__15735\,
            in3 => \N__10082\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22000\,
            ce => 'H',
            sr => \N__22298\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_15_LC_3_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12469\,
            in1 => \N__12349\,
            in2 => \N__15736\,
            in3 => \N__10061\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22000\,
            ce => 'H',
            sr => \N__22298\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_14_LC_3_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12345\,
            in1 => \N__15715\,
            in2 => \N__12496\,
            in3 => \N__10040\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22000\,
            ce => 'H',
            sr => \N__22298\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_12_LC_3_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12344\,
            in1 => \N__15714\,
            in2 => \N__12495\,
            in3 => \N__10019\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22000\,
            ce => 'H',
            sr => \N__22298\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_19_LC_3_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__12293\,
            in1 => \N__15703\,
            in2 => \N__12464\,
            in3 => \N__10238\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21995\,
            ce => 'H',
            sr => \N__22301\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_17_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12414\,
            in1 => \N__12294\,
            in2 => \N__15731\,
            in3 => \N__10217\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21995\,
            ce => 'H',
            sr => \N__22301\
        );

    \phase_controller_slave.stoper_hc.accumulated_time_18_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__12415\,
            in1 => \N__12295\,
            in2 => \N__15732\,
            in3 => \N__10196\,
            lcout => \phase_controller_slave.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21995\,
            ce => 'H',
            sr => \N__22301\
        );

    \phase_controller_slave.stoper_hc.stoper_state_0_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__12416\,
            in1 => \N__12296\,
            in2 => \N__15733\,
            in3 => \N__18060\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21992\,
            ce => \N__21289\,
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_1_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__18061\,
            in1 => \N__15710\,
            in2 => \N__12341\,
            in3 => \N__12417\,
            lcout => \phase_controller_slave.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21992\,
            ce => \N__21289\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_12_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11321\,
            in1 => \N__20939\,
            in2 => \_gnd_net_\,
            in3 => \N__10589\,
            lcout => measured_delay_tr_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22040\,
            ce => \N__11281\,
            sr => \N__22241\
        );

    \delay_measurement_inst.delay_tr_reg_esr_10_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__20937\,
            in1 => \N__11322\,
            in2 => \_gnd_net_\,
            in3 => \N__10628\,
            lcout => measured_delay_tr_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22040\,
            ce => \N__11281\,
            sr => \N__22241\
        );

    \delay_measurement_inst.delay_tr_reg_esr_11_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11320\,
            in1 => \N__20938\,
            in2 => \_gnd_net_\,
            in3 => \N__10610\,
            lcout => measured_delay_tr_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22040\,
            ce => \N__11281\,
            sr => \N__22241\
        );

    \delay_measurement_inst.tr_state_RNI5KUTL_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__11060\,
            in1 => \N__10262\,
            in2 => \N__20873\,
            in3 => \N__10175\,
            lcout => \delay_measurement_inst.N_81_i\,
            ltout => \delay_measurement_inst.N_81_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_RNICTS5M_0_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10160\,
            in3 => \N__22335\,
            lcout => \delay_measurement_inst.N_81_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA9RL2_15_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__10519\,
            in2 => \_gnd_net_\,
            in3 => \N__10455\,
            lcout => \delay_measurement_inst.N_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110001"
        )
    port map (
            in0 => \N__10562\,
            in1 => \N__10520\,
            in2 => \N__10456\,
            in3 => \N__11377\,
            lcout => \delay_measurement_inst.N_197_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_15_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__13677\,
            in1 => \N__13719\,
            in2 => \N__13784\,
            in3 => \N__13640\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_0_6_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13008\,
            in1 => \N__12603\,
            in2 => \N__12987\,
            in3 => \N__12873\,
            lcout => \phase_controller_inst1.stoper_tr.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011100"
        )
    port map (
            in0 => \N__11378\,
            in1 => \N__20936\,
            in2 => \N__10457\,
            in3 => \N__10244\,
            lcout => \delay_measurement_inst.N_165\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBIVI2_3_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10564\,
            in1 => \N__10448\,
            in2 => \N__10411\,
            in3 => \N__10424\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAFV93_7_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10271\,
            in1 => \N__10303\,
            in2 => \N__10265\,
            in3 => \N__10330\,
            lcout => \delay_measurement_inst.un1_tr_state_1_i_0_a2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10588\,
            in1 => \N__10609\,
            in2 => \N__11303\,
            in3 => \N__10624\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10\,
            ltout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__11094\,
            in1 => \N__10518\,
            in2 => \N__10247\,
            in3 => \N__10565\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__10477\,
            in1 => \N__11427\,
            in2 => \N__11405\,
            in3 => \N__11449\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_0_16_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11448\,
            in1 => \N__11400\,
            in2 => \N__11429\,
            in3 => \N__10476\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10381\,
            in2 => \_gnd_net_\,
            in3 => \N__10960\,
            lcout => \delay_measurement_inst.delay_tr_timer.un1_tr_state_1_i_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11242\,
            in2 => \N__11188\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11209\,
            in2 => \N__11164\,
            in3 => \N__10388\,
            lcout => \delay_measurement_inst.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11139\,
            in2 => \N__11189\,
            in3 => \N__10370\,
            lcout => \delay_measurement_inst.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11625\,
            in2 => \N__11165\,
            in3 => \N__10337\,
            lcout => \delay_measurement_inst.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11140\,
            in2 => \N__11608\,
            in3 => \N__10313\,
            lcout => \delay_measurement_inst.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11626\,
            in2 => \N__11584\,
            in3 => \N__10286\,
            lcout => \delay_measurement_inst.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11559\,
            in2 => \N__11609\,
            in3 => \N__10631\,
            lcout => \delay_measurement_inst.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11540\,
            in2 => \N__11585\,
            in3 => \N__10613\,
            lcout => \delay_measurement_inst.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__22032\,
            ce => \N__10726\,
            sr => \N__22255\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11561\,
            in2 => \N__11515\,
            in3 => \N__10592\,
            lcout => \delay_measurement_inst.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11539\,
            in2 => \N__11491\,
            in3 => \N__10571\,
            lcout => \delay_measurement_inst.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11466\,
            in2 => \N__11516\,
            in3 => \N__10568\,
            lcout => \delay_measurement_inst.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11820\,
            in2 => \N__11492\,
            in3 => \N__10532\,
            lcout => \delay_measurement_inst.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11467\,
            in2 => \N__11803\,
            in3 => \N__10484\,
            lcout => \delay_measurement_inst.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11821\,
            in2 => \N__11779\,
            in3 => \N__10460\,
            lcout => \delay_measurement_inst.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11756\,
            in2 => \N__11804\,
            in3 => \N__10694\,
            lcout => \delay_measurement_inst.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11732\,
            in2 => \N__11780\,
            in3 => \N__10691\,
            lcout => \delay_measurement_inst.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__22027\,
            ce => \N__10725\,
            sr => \N__22262\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11755\,
            in2 => \N__11707\,
            in3 => \N__10688\,
            lcout => \delay_measurement_inst.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_4_17_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_4_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11731\,
            in2 => \N__11683\,
            in3 => \N__10679\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11658\,
            in2 => \N__11708\,
            in3 => \N__10670\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_4_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11640\,
            in2 => \N__11684\,
            in3 => \N__10661\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11659\,
            in2 => \N__12133\,
            in3 => \N__10652\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_4_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11641\,
            in2 => \N__12109\,
            in3 => \N__10643\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12086\,
            in2 => \N__12134\,
            in3 => \N__10634\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_4_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12062\,
            in2 => \N__12110\,
            in3 => \N__10772\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__22023\,
            ce => \N__10724\,
            sr => \N__22271\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12085\,
            in2 => \N__12037\,
            in3 => \N__10763\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_4_18_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__22019\,
            ce => \N__10723\,
            sr => \N__22275\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12061\,
            in2 => \N__12013\,
            in3 => \N__10754\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__22019\,
            ce => \N__10723\,
            sr => \N__22275\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11989\,
            in2 => \N__12038\,
            in3 => \N__10745\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__22019\,
            ce => \N__10723\,
            sr => \N__22275\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11851\,
            in2 => \N__12014\,
            in3 => \N__10733\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__22019\,
            ce => \N__10723\,
            sr => \N__22275\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_4_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10730\,
            lcout => \delay_measurement_inst.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22019\,
            ce => \N__10723\,
            sr => \N__22275\
        );

    \phase_controller_slave.stoper_hc.target_time_5_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15353\,
            in1 => \N__14731\,
            in2 => \_gnd_net_\,
            in3 => \N__15455\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_3_LC_4_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__15580\,
            in1 => \N__13591\,
            in2 => \N__15920\,
            in3 => \N__14665\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_7_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15354\,
            in1 => \N__16148\,
            in2 => \_gnd_net_\,
            in3 => \N__15456\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_2_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15453\,
            in1 => \N__13589\,
            in2 => \N__16106\,
            in3 => \N__15356\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_1_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__13590\,
            in1 => \N__15916\,
            in2 => \N__14222\,
            in3 => \N__15579\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_0_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15452\,
            in1 => \N__13588\,
            in2 => \N__14129\,
            in3 => \N__15355\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_timeZ0Z_6_LC_4_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__14569\,
            in1 => \N__15915\,
            in2 => \_gnd_net_\,
            in3 => \N__15578\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_4_LC_4_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15454\,
            in1 => \N__15352\,
            in2 => \_gnd_net_\,
            in3 => \N__14264\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22014\,
            ce => \N__12245\,
            sr => \N__22279\
        );

    \phase_controller_slave.stoper_hc.target_time_12_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15331\,
            in1 => \N__16013\,
            in2 => \_gnd_net_\,
            in3 => \N__15436\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22008\,
            ce => \N__12241\,
            sr => \N__22285\
        );

    \phase_controller_slave.stoper_hc.target_time_10_LC_4_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15329\,
            in1 => \N__15965\,
            in2 => \_gnd_net_\,
            in3 => \N__15434\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22008\,
            ce => \N__12241\,
            sr => \N__22285\
        );

    \phase_controller_slave.stoper_hc.target_time_13_LC_4_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15437\,
            in1 => \N__15332\,
            in2 => \_gnd_net_\,
            in3 => \N__14510\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22008\,
            ce => \N__12241\,
            sr => \N__22285\
        );

    \phase_controller_slave.stoper_hc.target_time_11_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15435\,
            in1 => \N__15330\,
            in2 => \_gnd_net_\,
            in3 => \N__15785\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22008\,
            ce => \N__12241\,
            sr => \N__22285\
        );

    \phase_controller_slave.stoper_hc.target_time_8_LC_4_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__16059\,
            in1 => \_gnd_net_\,
            in2 => \N__15357\,
            in3 => \N__15439\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22008\,
            ce => \N__12241\,
            sr => \N__22285\
        );

    \phase_controller_slave.stoper_hc.target_time_15_LC_4_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15438\,
            in1 => \N__15333\,
            in2 => \_gnd_net_\,
            in3 => \N__14398\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22008\,
            ce => \N__12241\,
            sr => \N__22285\
        );

    \phase_controller_slave.stoper_hc.target_time_14_LC_4_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__15895\,
            in1 => \N__14830\,
            in2 => \_gnd_net_\,
            in3 => \N__15553\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22001\,
            ce => \N__12240\,
            sr => \N__22290\
        );

    \phase_controller_slave.stoper_hc.target_time_9_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__15554\,
            in1 => \N__15896\,
            in2 => \_gnd_net_\,
            in3 => \N__16195\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22001\,
            ce => \N__12240\,
            sr => \N__22290\
        );

    \phase_controller_slave.stoper_hc.target_time_19_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__14457\,
            in1 => \N__15892\,
            in2 => \_gnd_net_\,
            in3 => \N__15533\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21996\,
            ce => \N__12239\,
            sr => \N__22294\
        );

    \phase_controller_slave.stoper_hc.target_time_18_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__15532\,
            in1 => \_gnd_net_\,
            in2 => \N__15906\,
            in3 => \N__14338\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21996\,
            ce => \N__12239\,
            sr => \N__22294\
        );

    \phase_controller_slave.stoper_hc.target_time_16_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__14875\,
            in1 => \N__15885\,
            in2 => \_gnd_net_\,
            in3 => \N__15530\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21996\,
            ce => \N__12239\,
            sr => \N__22294\
        );

    \phase_controller_slave.stoper_hc.target_time_17_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001010"
        )
    port map (
            in0 => \N__15531\,
            in1 => \_gnd_net_\,
            in2 => \N__15905\,
            in3 => \N__14616\,
            lcout => \phase_controller_slave.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21996\,
            ce => \N__12239\,
            sr => \N__22294\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_7_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14876\,
            in1 => \N__14507\,
            in2 => \N__14570\,
            in3 => \N__15959\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_8_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14339\,
            in1 => \N__14722\,
            in2 => \N__14459\,
            in3 => \N__14262\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_10_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16139\,
            in1 => \N__16006\,
            in2 => \N__16061\,
            in3 => \N__15778\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_15_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12644\,
            in1 => \N__18735\,
            in2 => \N__10949\,
            in3 => \N__18691\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10946\,
            in1 => \N__10940\,
            in2 => \N__10934\,
            in3 => \N__12668\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlt31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNIDEUE_0_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12396\,
            in2 => \_gnd_net_\,
            in3 => \N__12279\,
            lcout => \phase_controller_slave.stoper_hc.time_passed11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D1_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MAX_D2_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10919\,
            lcout => \il_max_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21485\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_6_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000101"
        )
    port map (
            in0 => \N__12957\,
            in1 => \N__12566\,
            in2 => \N__20027\,
            in3 => \N__12535\,
            lcout => \phase_controller_inst1.stoper_tr.N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_3_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13676\,
            in1 => \N__13718\,
            in2 => \N__13769\,
            in3 => \N__13644\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4_3_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12956\,
            in1 => \N__12739\,
            in2 => \N__20026\,
            in3 => \N__12843\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_4Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6_3_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__12822\,
            in1 => \N__11111\,
            in2 => \N__11123\,
            in3 => \N__11120\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_6Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f0_0_0_a2_3_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12567\,
            in2 => \N__11114\,
            in3 => \N__12537\,
            lcout => \phase_controller_inst1.stoper_tr.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0_6_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12778\,
            in2 => \_gnd_net_\,
            in3 => \N__13179\,
            lcout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6\,
            ltout => \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a2_1_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_0_a3_0_6_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20014\,
            in1 => \N__12823\,
            in2 => \N__11105\,
            in3 => \N__12536\,
            lcout => \phase_controller_inst1.stoper_tr.N_92\,
            ltout => \phase_controller_inst1.stoper_tr.N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_i_0_o2_2_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__20071\,
            in1 => \_gnd_net_\,
            in2 => \N__11102\,
            in3 => \N__13118\,
            lcout => \phase_controller_inst1.stoper_tr.N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_reg_esr_9_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__20947\,
            in1 => \N__11324\,
            in2 => \N__11099\,
            in3 => \N__11071\,
            lcout => measured_delay_tr_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22033\,
            ce => \N__11282\,
            sr => \N__22243\
        );

    \delay_measurement_inst.delay_tr_reg_esr_4_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__11072\,
            in1 => \N__11035\,
            in2 => \N__11000\,
            in3 => \N__10961\,
            lcout => measured_delay_tr_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22033\,
            ce => \N__11282\,
            sr => \N__22243\
        );

    \delay_measurement_inst.delay_tr_reg_esr_18_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__20945\,
            in1 => \N__11450\,
            in2 => \_gnd_net_\,
            in3 => \N__11380\,
            lcout => measured_delay_tr_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22033\,
            ce => \N__11282\,
            sr => \N__22243\
        );

    \delay_measurement_inst.delay_tr_reg_esr_19_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__11381\,
            in1 => \N__20946\,
            in2 => \_gnd_net_\,
            in3 => \N__11428\,
            lcout => measured_delay_tr_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22033\,
            ce => \N__11282\,
            sr => \N__22243\
        );

    \delay_measurement_inst.delay_tr_reg_esr_17_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__20944\,
            in1 => \N__11404\,
            in2 => \_gnd_net_\,
            in3 => \N__11379\,
            lcout => measured_delay_tr_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22033\,
            ce => \N__11282\,
            sr => \N__22243\
        );

    \delay_measurement_inst.delay_tr_reg_esr_13_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__11323\,
            in1 => \N__20943\,
            in2 => \_gnd_net_\,
            in3 => \N__11302\,
            lcout => measured_delay_tr_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22033\,
            ce => \N__11282\,
            sr => \N__22243\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11972\,
            in1 => \N__11235\,
            in2 => \_gnd_net_\,
            in3 => \N__11219\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11968\,
            in1 => \N__11208\,
            in2 => \_gnd_net_\,
            in3 => \N__11192\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11973\,
            in1 => \N__11187\,
            in2 => \_gnd_net_\,
            in3 => \N__11168\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11969\,
            in1 => \N__11163\,
            in2 => \_gnd_net_\,
            in3 => \N__11144\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11974\,
            in1 => \N__11141\,
            in2 => \_gnd_net_\,
            in3 => \N__11126\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11970\,
            in1 => \N__11627\,
            in2 => \_gnd_net_\,
            in3 => \N__11612\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11975\,
            in1 => \N__11607\,
            in2 => \_gnd_net_\,
            in3 => \N__11588\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11971\,
            in1 => \N__11583\,
            in2 => \_gnd_net_\,
            in3 => \N__11564\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__22028\,
            ce => \N__11837\,
            sr => \N__22249\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11949\,
            in1 => \N__11560\,
            in2 => \_gnd_net_\,
            in3 => \N__11543\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11953\,
            in1 => \N__11538\,
            in2 => \_gnd_net_\,
            in3 => \N__11519\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11946\,
            in1 => \N__11514\,
            in2 => \_gnd_net_\,
            in3 => \N__11495\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11950\,
            in1 => \N__11490\,
            in2 => \_gnd_net_\,
            in3 => \N__11471\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11947\,
            in1 => \N__11468\,
            in2 => \_gnd_net_\,
            in3 => \N__11453\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11951\,
            in1 => \N__11822\,
            in2 => \_gnd_net_\,
            in3 => \N__11807\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11948\,
            in1 => \N__11802\,
            in2 => \_gnd_net_\,
            in3 => \N__11783\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11952\,
            in1 => \N__11778\,
            in2 => \_gnd_net_\,
            in3 => \N__11759\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__22024\,
            ce => \N__11838\,
            sr => \N__22256\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11954\,
            in1 => \N__11754\,
            in2 => \_gnd_net_\,
            in3 => \N__11735\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_5_17_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11958\,
            in1 => \N__11730\,
            in2 => \_gnd_net_\,
            in3 => \N__11711\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11955\,
            in1 => \N__11706\,
            in2 => \_gnd_net_\,
            in3 => \N__11687\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11959\,
            in1 => \N__11682\,
            in2 => \_gnd_net_\,
            in3 => \N__11663\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11956\,
            in1 => \N__11660\,
            in2 => \_gnd_net_\,
            in3 => \N__11645\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11960\,
            in1 => \N__11642\,
            in2 => \_gnd_net_\,
            in3 => \N__12137\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11957\,
            in1 => \N__12132\,
            in2 => \_gnd_net_\,
            in3 => \N__12113\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11961\,
            in1 => \N__12108\,
            in2 => \_gnd_net_\,
            in3 => \N__12089\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__22020\,
            ce => \N__11839\,
            sr => \N__22263\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11962\,
            in1 => \N__12084\,
            in2 => \_gnd_net_\,
            in3 => \N__12065\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_5_18_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__22015\,
            ce => \N__11840\,
            sr => \N__22272\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11966\,
            in1 => \N__12060\,
            in2 => \_gnd_net_\,
            in3 => \N__12041\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__22015\,
            ce => \N__11840\,
            sr => \N__22272\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11963\,
            in1 => \N__12036\,
            in2 => \_gnd_net_\,
            in3 => \N__12017\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__22015\,
            ce => \N__11840\,
            sr => \N__22272\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11967\,
            in1 => \N__12012\,
            in2 => \_gnd_net_\,
            in3 => \N__11993\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__22015\,
            ce => \N__11840\,
            sr => \N__22272\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11964\,
            in1 => \N__11990\,
            in2 => \_gnd_net_\,
            in3 => \N__11978\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__22015\,
            ce => \N__11840\,
            sr => \N__22272\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11852\,
            in1 => \N__11965\,
            in2 => \_gnd_net_\,
            in3 => \N__11855\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22015\,
            ce => \N__11840\,
            sr => \N__22272\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15450\,
            in1 => \N__15350\,
            in2 => \_gnd_net_\,
            in3 => \N__14732\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22009\,
            ce => \N__18499\,
            sr => \N__22276\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15351\,
            in1 => \N__16147\,
            in2 => \_gnd_net_\,
            in3 => \N__15451\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22009\,
            ce => \N__18499\,
            sr => \N__22276\
        );

    \phase_controller_inst1.stoper_hc.target_timeZ0Z_6_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__14565\,
            in1 => \N__15907\,
            in2 => \_gnd_net_\,
            in3 => \N__15576\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22009\,
            ce => \N__18499\,
            sr => \N__22276\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15349\,
            in1 => \N__14263\,
            in2 => \_gnd_net_\,
            in3 => \N__15449\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22009\,
            ce => \N__18499\,
            sr => \N__22276\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15412\,
            in1 => \N__15310\,
            in2 => \_gnd_net_\,
            in3 => \N__14399\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22002\,
            ce => \N__18500\,
            sr => \N__22280\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15309\,
            in1 => \N__15411\,
            in2 => \_gnd_net_\,
            in3 => \N__14509\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22002\,
            ce => \N__18500\,
            sr => \N__22280\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_d_0_LC_5_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110110011"
        )
    port map (
            in0 => \N__12515\,
            in1 => \N__12184\,
            in2 => \N__12146\,
            in3 => \N__12161\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto31_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.time_passed_RNO_0_LC_5_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15665\,
            in1 => \N__12465\,
            in2 => \_gnd_net_\,
            in3 => \N__12342\,
            lcout => \phase_controller_slave.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un3_start_0_a0_0_LC_5_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18740\,
            in1 => \N__18710\,
            in2 => \N__12662\,
            in3 => \N__15894\,
            lcout => \phase_controller_inst1.stoper_hc.un3_start_0_a0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m3_e_1_LC_5_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__15893\,
            in1 => \N__14393\,
            in2 => \_gnd_net_\,
            in3 => \N__14829\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m3_eZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m3_0_1_LC_5_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16009\,
            in1 => \N__15784\,
            in2 => \N__14508\,
            in3 => \N__15961\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_a0_1_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15884\,
            in1 => \N__14831\,
            in2 => \_gnd_net_\,
            in3 => \N__12514\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto31_a0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto19_2_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14333\,
            in1 => \N__14615\,
            in2 => \N__14458\,
            in3 => \N__14874\,
            lcout => phase_controller_inst1_stoper_hc_un1_startlto19_2,
            ltout => \phase_controller_inst1_stoper_hc_un1_startlto19_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_1_RNIQA9D_15_LC_5_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15882\,
            in2 => \N__12503\,
            in3 => \N__14392\,
            lcout => \d_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_hc.stoper_state_RNI10KL_0_LC_5_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__15698\,
            in1 => \N__12466\,
            in2 => \_gnd_net_\,
            in3 => \N__12343\,
            lcout => \phase_controller_slave.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_a2_LC_5_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__12655\,
            in1 => \N__18736\,
            in2 => \N__18709\,
            in3 => \N__15883\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_startlto31_aZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto31_1_LC_5_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__12194\,
            in1 => \N__12160\,
            in2 => \N__12188\,
            in3 => \N__12185\,
            lcout => \phase_controller_inst1.stoper_hc.un1_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m3_0_2_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__16138\,
            in1 => \N__16045\,
            in2 => \N__16196\,
            in3 => \N__12173\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_m3_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m3_0_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__14554\,
            in1 => \N__16194\,
            in2 => \N__12164\,
            in3 => \N__12677\,
            lcout => \phase_controller_inst1.stoper_hc.un1_N_6_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_3_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14252\,
            in1 => \N__14651\,
            in2 => \N__14730\,
            in3 => \N__14121\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_m2_e_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__14206\,
            in1 => \_gnd_net_\,
            in2 => \N__12680\,
            in3 => \N__16094\,
            lcout => \phase_controller_inst1.stoper_hc.un1_m2_eZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_6_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__16190\,
            in1 => \N__14684\,
            in2 => \_gnd_net_\,
            in3 => \N__14617\,
            lcout => OPEN,
            ltout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_11_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__14207\,
            in1 => \N__14652\,
            in2 => \N__12671\,
            in3 => \N__16095\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_startlto30_2_0_0_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14149\,
            in1 => \N__14170\,
            in2 => \_gnd_net_\,
            in3 => \N__14683\,
            lcout => \phase_controller_inst1.stoper_hc.un1_startlto30_2_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_9_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14171\,
            in1 => \N__14828\,
            in2 => \N__14397\,
            in3 => \N__14150\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_5_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12923\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12610\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22034\,
            ce => \N__19944\,
            sr => \N__22233\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011110011"
        )
    port map (
            in0 => \N__20032\,
            in1 => \N__12926\,
            in2 => \N__12587\,
            in3 => \N__12548\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22034\,
            ce => \N__19944\,
            sr => \N__22233\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13015\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22034\,
            ce => \N__19944\,
            sr => \N__22233\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12925\,
            in2 => \_gnd_net_\,
            in3 => \N__12995\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22034\,
            ce => \N__19944\,
            sr => \N__22233\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__20031\,
            in2 => \_gnd_net_\,
            in3 => \N__12962\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22034\,
            ce => \N__19944\,
            sr => \N__22233\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12922\,
            in2 => \_gnd_net_\,
            in3 => \N__12880\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22034\,
            ce => \N__19944\,
            sr => \N__22233\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__13138\,
            in1 => \N__20118\,
            in2 => \N__13234\,
            in3 => \N__12856\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12827\,
            in1 => \N__20116\,
            in2 => \_gnd_net_\,
            in3 => \N__13136\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__13137\,
            in1 => \N__20117\,
            in2 => \_gnd_net_\,
            in3 => \N__12782\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__20119\,
            in1 => \N__12743\,
            in2 => \N__13233\,
            in3 => \N__13139\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__12719\,
            in1 => \N__13289\,
            in2 => \N__12701\,
            in3 => \N__13264\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__13263\,
            in1 => \N__13337\,
            in2 => \N__13301\,
            in3 => \N__13358\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__13336\,
            in1 => \N__13293\,
            in2 => \_gnd_net_\,
            in3 => \N__13265\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000000110001"
        )
    port map (
            in0 => \N__20120\,
            in1 => \N__13224\,
            in2 => \N__13187\,
            in3 => \N__13140\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22029\,
            ce => \N__19949\,
            sr => \N__22237\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13100\,
            in2 => \N__13094\,
            in3 => \N__17067\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13085\,
            in2 => \N__13076\,
            in3 => \N__17035\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13067\,
            in2 => \N__13061\,
            in3 => \N__17014\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13052\,
            in2 => \N__13046\,
            in3 => \N__16981\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16960\,
            in1 => \N__13037\,
            in2 => \N__13028\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13487\,
            in2 => \N__13481\,
            in3 => \N__16939\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17290\,
            in1 => \N__13472\,
            in2 => \N__13466\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17269\,
            in1 => \N__13457\,
            in2 => \N__13448\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13439\,
            in2 => \N__13430\,
            in3 => \N__17248\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13421\,
            in2 => \N__13412\,
            in3 => \N__17227\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13403\,
            in2 => \N__13394\,
            in3 => \N__17203\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13385\,
            in2 => \N__13376\,
            in3 => \N__17183\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13367\,
            in2 => \N__13565\,
            in3 => \N__17155\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13556\,
            in2 => \N__13547\,
            in3 => \N__17131\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19961\,
            in2 => \N__13538\,
            in3 => \N__17668\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13616\,
            in2 => \N__13529\,
            in3 => \N__17644\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13697\,
            in2 => \N__13520\,
            in3 => \N__17623\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13658\,
            in2 => \N__13511\,
            in3 => \N__17602\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13739\,
            in2 => \N__13502\,
            in3 => \N__17581\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13493\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13490\,
            in3 => \N__19734\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_RNII60D_0_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__15237\,
            in1 => \_gnd_net_\,
            in2 => \N__15008\,
            in3 => \N__19789\,
            lcout => \phase_controller_slave.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13782\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22010\,
            ce => \N__19929\,
            sr => \N__22250\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13733\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22010\,
            ce => \N__19929\,
            sr => \N__22250\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13691\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22010\,
            ce => \N__19929\,
            sr => \N__22250\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13652\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22010\,
            ce => \N__19929\,
            sr => \N__22250\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__15903\,
            in1 => \N__13606\,
            in2 => \N__14221\,
            in3 => \N__15586\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22003\,
            ce => \N__18487\,
            sr => \N__22257\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__15904\,
            in1 => \N__15587\,
            in2 => \N__14666\,
            in3 => \N__13607\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22003\,
            ce => \N__18487\,
            sr => \N__22257\
        );

    \phase_controller_inst1.stoper_hc.target_time_0_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13604\,
            in1 => \N__14122\,
            in2 => \N__15373\,
            in3 => \N__15466\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22003\,
            ce => \N__18487\,
            sr => \N__22257\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13605\,
            in1 => \N__16102\,
            in2 => \N__15374\,
            in3 => \N__15467\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22003\,
            ce => \N__18487\,
            sr => \N__22257\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13949\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13940\,
            in2 => \N__13934\,
            in3 => \N__18414\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13925\,
            in2 => \N__13919\,
            in3 => \N__17311\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13910\,
            in2 => \N__13904\,
            in3 => \N__17866\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13895\,
            in2 => \N__13886\,
            in3 => \N__17827\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13877\,
            in2 => \N__13868\,
            in3 => \N__17806\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17785\,
            in1 => \N__13859\,
            in2 => \N__13850\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17764\,
            in1 => \N__13841\,
            in2 => \N__13832\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15473\,
            in2 => \N__14042\,
            in3 => \N__17737\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15497\,
            in2 => \N__14033\,
            in3 => \N__17710\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15491\,
            in2 => \N__14024\,
            in3 => \N__17689\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15482\,
            in2 => \N__14015\,
            in3 => \N__18031\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15269\,
            in2 => \N__14006\,
            in3 => \N__18010\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13997\,
            in2 => \N__13988\,
            in3 => \N__17989\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14279\,
            in2 => \N__13979\,
            in3 => \N__17968\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17947\,
            in1 => \N__13970\,
            in2 => \N__13958\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17927\,
            in1 => \N__14048\,
            in2 => \N__14090\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_16\,
            ltout => OPEN,
            carryin => \bfn_7_21_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14288\,
            in2 => \N__14081\,
            in3 => \N__17902\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_17\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14297\,
            in2 => \N__14072\,
            in3 => \N__17878\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18520\,
            in1 => \N__14270\,
            in2 => \N__14063\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14054\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18438\,
            in2 => \_gnd_net_\,
            in3 => \N__18387\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18267\,
            in2 => \_gnd_net_\,
            in3 => \N__18163\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed11\,
            ltout => \phase_controller_inst1.stoper_hc.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14051\,
            in3 => \N__18388\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__15873\,
            in1 => \N__14873\,
            in2 => \_gnd_net_\,
            in3 => \N__15559\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21985\,
            ce => \N__18491\,
            sr => \N__22281\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__15561\,
            in1 => \N__15875\,
            in2 => \_gnd_net_\,
            in3 => \N__14337\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21985\,
            ce => \N__18491\,
            sr => \N__22281\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__15874\,
            in1 => \N__14614\,
            in2 => \_gnd_net_\,
            in3 => \N__15560\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21985\,
            ce => \N__18491\,
            sr => \N__22281\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__15872\,
            in1 => \N__14824\,
            in2 => \_gnd_net_\,
            in3 => \N__15558\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21985\,
            ce => \N__18491\,
            sr => \N__22281\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_7_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__15562\,
            in1 => \N__15876\,
            in2 => \_gnd_net_\,
            in3 => \N__14449\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21985\,
            ce => \N__18491\,
            sr => \N__22281\
        );

    \delay_measurement_inst.delay_hc_reg_4_LC_7_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__14251\,
            in1 => \N__19104\,
            in2 => \N__16277\,
            in3 => \N__18611\,
            lcout => measured_delay_hc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_1_LC_7_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__19102\,
            in1 => \N__18914\,
            in2 => \N__14214\,
            in3 => \N__18990\,
            lcout => measured_delay_hc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_22_LC_7_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18993\,
            in1 => \N__14169\,
            in2 => \_gnd_net_\,
            in3 => \N__19101\,
            lcout => measured_delay_hc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_21_LC_7_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19100\,
            in1 => \N__14148\,
            in2 => \_gnd_net_\,
            in3 => \N__18992\,
            lcout => measured_delay_hc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_0_LC_7_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14120\,
            in1 => \N__19098\,
            in2 => \_gnd_net_\,
            in3 => \N__18610\,
            lcout => measured_delay_hc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_5_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__19105\,
            in1 => \N__16606\,
            in2 => \N__14729\,
            in3 => \N__18995\,
            lcout => measured_delay_hc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_20_LC_7_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18991\,
            in1 => \N__14682\,
            in2 => \_gnd_net_\,
            in3 => \N__19099\,
            lcout => measured_delay_hc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_3_LC_7_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__19103\,
            in1 => \N__14650\,
            in2 => \N__16304\,
            in3 => \N__18994\,
            lcout => measured_delay_hc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21982\,
            ce => 'H',
            sr => \N__22286\
        );

    \delay_measurement_inst.delay_hc_reg_17_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011111010"
        )
    port map (
            in0 => \N__18603\,
            in1 => \N__16721\,
            in2 => \N__14618\,
            in3 => \N__19110\,
            lcout => measured_delay_hc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_6_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__19113\,
            in1 => \N__16577\,
            in2 => \N__14558\,
            in3 => \N__18606\,
            lcout => measured_delay_hc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_13_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__16400\,
            in1 => \N__19106\,
            in2 => \N__14497\,
            in3 => \N__18983\,
            lcout => measured_delay_hc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_19_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__19112\,
            in1 => \N__16667\,
            in2 => \N__14450\,
            in3 => \N__18605\,
            lcout => measured_delay_hc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_15_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000000000"
        )
    port map (
            in0 => \N__16798\,
            in1 => \N__19108\,
            in2 => \N__14385\,
            in3 => \N__18984\,
            lcout => measured_delay_hc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_18_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__19111\,
            in1 => \N__16694\,
            in2 => \N__14332\,
            in3 => \N__18604\,
            lcout => measured_delay_hc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_16_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__14863\,
            in2 => \N__16751\,
            in3 => \N__19109\,
            lcout => measured_delay_hc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_reg_14_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__19107\,
            in1 => \N__14814\,
            in2 => \N__16838\,
            in3 => \N__18601\,
            lcout => measured_delay_hc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21979\,
            ce => 'H',
            sr => \N__22291\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINAE19_14_LC_7_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__16322\,
            in1 => \N__14774\,
            in2 => \N__14762\,
            in3 => \N__14741\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_13_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16596\,
            in1 => \N__16263\,
            in2 => \N__16746\,
            in3 => \N__16392\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILU0I2_19_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16662\,
            in1 => \N__16573\,
            in2 => \N__14777\,
            in3 => \N__14768\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI537G_17_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16683\,
            in2 => \_gnd_net_\,
            in3 => \N__16710\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILLI01_20_LC_7_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16619\,
            in1 => \N__17083\,
            in2 => \N__16919\,
            in3 => \N__16633\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_7_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14909\,
            in1 => \N__14750\,
            in2 => \N__16637\,
            in3 => \N__14903\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto30_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_7_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16886\,
            in1 => \N__16895\,
            in2 => \N__16877\,
            in3 => \N__16904\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC512_23_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14744\,
            in3 => \N__14902\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16915\,
            in2 => \_gnd_net_\,
            in3 => \N__16618\,
            lcout => \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_7_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16847\,
            in1 => \N__16856\,
            in2 => \N__17111\,
            in3 => \N__16865\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lt31_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D1_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14894\,
            lcout => \il_min_comp2_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__17543\,
            in1 => \N__17431\,
            in2 => \N__20846\,
            in3 => \N__17258\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17426\,
            in1 => \N__20825\,
            in2 => \N__17559\,
            in3 => \N__16949\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__17542\,
            in1 => \N__17430\,
            in2 => \N__20845\,
            in3 => \N__16970\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17428\,
            in1 => \N__20827\,
            in2 => \N__17561\,
            in3 => \N__17279\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__17541\,
            in1 => \N__17429\,
            in2 => \N__20844\,
            in3 => \N__17024\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17427\,
            in1 => \N__20826\,
            in2 => \N__17560\,
            in3 => \N__16928\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17425\,
            in1 => \N__20824\,
            in2 => \N__17558\,
            in3 => \N__16991\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22025\,
            ce => 'H',
            sr => \N__22234\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17403\,
            in1 => \N__17532\,
            in2 => \N__20840\,
            in3 => \N__17237\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__17525\,
            in1 => \N__20808\,
            in2 => \N__17216\,
            in3 => \N__17404\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17401\,
            in1 => \N__17530\,
            in2 => \N__20838\,
            in3 => \N__17165\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__17527\,
            in1 => \N__20810\,
            in2 => \N__17657\,
            in3 => \N__17406\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17400\,
            in1 => \N__17529\,
            in2 => \N__20837\,
            in3 => \N__17192\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100100000000"
        )
    port map (
            in0 => \N__17528\,
            in1 => \N__20811\,
            in2 => \N__17435\,
            in3 => \N__17633\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17402\,
            in1 => \N__17531\,
            in2 => \N__20839\,
            in3 => \N__17120\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__17526\,
            in1 => \N__20809\,
            in2 => \N__17144\,
            in3 => \N__17405\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22021\,
            ce => 'H',
            sr => \N__22238\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17394\,
            in1 => \N__20813\,
            in2 => \N__17556\,
            in3 => \N__17591\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22016\,
            ce => 'H',
            sr => \N__22239\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__17540\,
            in1 => \N__17397\,
            in2 => \N__20842\,
            in3 => \N__14927\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22016\,
            ce => 'H',
            sr => \N__22239\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__17395\,
            in1 => \N__20814\,
            in2 => \N__17557\,
            in3 => \N__17567\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22016\,
            ce => 'H',
            sr => \N__22239\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__17539\,
            in1 => \N__17396\,
            in2 => \N__20841\,
            in3 => \N__17612\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22016\,
            ce => 'H',
            sr => \N__22239\
        );

    \phase_controller_slave.stoper_tr.time_passed_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__20487\,
            in1 => \N__14960\,
            in2 => \N__14918\,
            in3 => \N__15122\,
            lcout => \phase_controller_slave.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22016\,
            ce => 'H',
            sr => \N__22239\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20779\,
            in1 => \N__17470\,
            in2 => \_gnd_net_\,
            in3 => \N__17371\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__19735\,
            in1 => \N__19706\,
            in2 => \_gnd_net_\,
            in3 => \N__17071\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17469\,
            in2 => \_gnd_net_\,
            in3 => \N__17370\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed11\,
            ltout => \phase_controller_inst1.stoper_tr.time_passed11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14921\,
            in3 => \N__19705\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.time_passed_RNO_0_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__19790\,
            in1 => \N__14997\,
            in2 => \_gnd_net_\,
            in3 => \N__15238\,
            lcout => \phase_controller_slave.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__17372\,
            in1 => \_gnd_net_\,
            in2 => \N__17508\,
            in3 => \N__20780\,
            lcout => \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.stoper_tr.stoper_state_1_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__15001\,
            in1 => \N__15258\,
            in2 => \N__19873\,
            in3 => \N__15118\,
            lcout => \phase_controller_slave.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22004\,
            ce => \N__21331\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_1_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001100100"
        )
    port map (
            in0 => \N__17506\,
            in1 => \N__17399\,
            in2 => \N__20843\,
            in3 => \N__19713\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22004\,
            ce => \N__21331\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18232\,
            in1 => \N__20634\,
            in2 => \N__18350\,
            in3 => \N__17753\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => 'H',
            sr => \N__22251\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18337\,
            in1 => \N__18235\,
            in2 => \N__20657\,
            in3 => \N__17774\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => 'H',
            sr => \N__22251\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18336\,
            in1 => \N__18234\,
            in2 => \N__20656\,
            in3 => \N__17795\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => 'H',
            sr => \N__22251\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18231\,
            in1 => \N__20633\,
            in2 => \N__18349\,
            in3 => \N__17816\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => 'H',
            sr => \N__22251\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18335\,
            in1 => \N__18233\,
            in2 => \N__20655\,
            in3 => \N__17300\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => 'H',
            sr => \N__22251\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18230\,
            in1 => \N__20632\,
            in2 => \N__18348\,
            in3 => \N__17837\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21997\,
            ce => 'H',
            sr => \N__22251\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18328\,
            in1 => \N__18227\,
            in2 => \N__20646\,
            in3 => \N__17957\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18223\,
            in1 => \N__18332\,
            in2 => \N__20652\,
            in3 => \N__18020\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18329\,
            in1 => \N__18228\,
            in2 => \N__20647\,
            in3 => \N__17936\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18225\,
            in1 => \N__18334\,
            in2 => \N__20654\,
            in3 => \N__17912\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18330\,
            in1 => \N__18229\,
            in2 => \N__20648\,
            in3 => \N__17699\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18222\,
            in1 => \N__18331\,
            in2 => \N__20651\,
            in3 => \N__17678\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18327\,
            in1 => \N__18226\,
            in2 => \N__20645\,
            in3 => \N__17999\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18224\,
            in1 => \N__18333\,
            in2 => \N__20653\,
            in3 => \N__17978\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21993\,
            ce => 'H',
            sr => \N__22258\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101100000000"
        )
    port map (
            in0 => \N__18218\,
            in1 => \N__18325\,
            in2 => \N__20650\,
            in3 => \N__18506\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__18324\,
            in1 => \N__20616\,
            in2 => \N__17726\,
            in3 => \N__18221\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__20403\,
            in1 => \N__18442\,
            in2 => \N__18134\,
            in3 => \N__18394\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010110000"
        )
    port map (
            in0 => \N__18217\,
            in1 => \N__20611\,
            in2 => \N__18533\,
            in3 => \N__18326\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__18322\,
            in1 => \N__20615\,
            in2 => \N__17891\,
            in3 => \N__18220\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_slave.start_timer_hc_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__15633\,
            in1 => \N__18356\,
            in2 => \N__20348\,
            in3 => \N__18125\,
            lcout => \phase_controller_slave.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110100000000"
        )
    port map (
            in0 => \N__18323\,
            in1 => \N__18219\,
            in2 => \N__20649\,
            in3 => \N__18362\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21990\,
            ce => 'H',
            sr => \N__22264\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__15871\,
            in1 => \N__16186\,
            in2 => \_gnd_net_\,
            in3 => \N__15577\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21986\,
            ce => \N__18492\,
            sr => \N__22273\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15358\,
            in1 => \N__15960\,
            in2 => \_gnd_net_\,
            in3 => \N__15462\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21986\,
            ce => \N__18492\,
            sr => \N__22273\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15463\,
            in1 => \N__15359\,
            in2 => \_gnd_net_\,
            in3 => \N__15779\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21986\,
            ce => \N__18492\,
            sr => \N__22273\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15361\,
            in1 => \N__16055\,
            in2 => \_gnd_net_\,
            in3 => \N__15465\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21986\,
            ce => \N__18492\,
            sr => \N__22273\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15464\,
            in1 => \N__15360\,
            in2 => \_gnd_net_\,
            in3 => \N__16007\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21986\,
            ce => \N__18492\,
            sr => \N__22273\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_0_LC_8_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__18316\,
            in1 => \N__18211\,
            in2 => \N__20644\,
            in3 => \N__18392\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21983\,
            ce => \N__21324\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_1_LC_8_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001010000"
        )
    port map (
            in0 => \N__18393\,
            in1 => \N__20595\,
            in2 => \N__18236\,
            in3 => \N__18317\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21983\,
            ce => \N__21324\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_9_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111011101"
        )
    port map (
            in0 => \N__18982\,
            in1 => \N__16185\,
            in2 => \N__16508\,
            in3 => \N__19097\,
            lcout => measured_delay_hc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_7_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__19095\,
            in1 => \N__18980\,
            in2 => \N__16146\,
            in3 => \N__16553\,
            lcout => measured_delay_hc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_2_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__18979\,
            in1 => \N__16093\,
            in2 => \N__18896\,
            in3 => \N__19094\,
            lcout => measured_delay_hc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_8_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__19096\,
            in1 => \N__16532\,
            in2 => \N__16060\,
            in3 => \N__18981\,
            lcout => measured_delay_hc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_12_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__18599\,
            in1 => \N__19093\,
            in2 => \N__16008\,
            in3 => \N__16427\,
            lcout => measured_delay_hc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_10_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__16472\,
            in1 => \N__15952\,
            in2 => \N__19118\,
            in3 => \N__18978\,
            lcout => measured_delay_hc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_31_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__18600\,
            in1 => \N__15838\,
            in2 => \_gnd_net_\,
            in3 => \N__19088\,
            lcout => measured_delay_hc_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_reg_11_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19092\,
            in1 => \N__18598\,
            in2 => \N__15783\,
            in3 => \N__16451\,
            lcout => measured_delay_hc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21980\,
            ce => 'H',
            sr => \N__22282\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_0_31_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__16216\,
            in1 => \N__16366\,
            in2 => \N__17096\,
            in3 => \N__16226\,
            lcout => \delay_measurement_inst.delay_hc_reg3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1_9_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16346\,
            in1 => \N__16503\,
            in2 => \_gnd_net_\,
            in3 => \N__16795\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5FBM1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI93LG1_14_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__16796\,
            in1 => \N__16832\,
            in2 => \_gnd_net_\,
            in3 => \N__16316\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIABFQE_14_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__16247\,
            in1 => \N__16202\,
            in2 => \N__16241\,
            in3 => \N__16238\,
            lcout => \delay_measurement_inst.un1_elapsed_time_hc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18907\,
            in1 => \N__16300\,
            in2 => \N__16607\,
            in3 => \N__18888\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FS83_4_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16270\,
            in1 => \N__16793\,
            in2 => \N__16232\,
            in3 => \N__16358\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_a0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9U7V4_9_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__16794\,
            in1 => \N__16507\,
            in2 => \N__16229\,
            in3 => \N__16345\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNINHL3C_31_LC_8_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__16367\,
            in1 => \N__17095\,
            in2 => \N__16220\,
            in3 => \N__16217\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto31_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2_6_LC_8_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16572\,
            in1 => \N__16344\,
            in2 => \N__16799\,
            in3 => \N__16357\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6\,
            ltout => \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5E0I2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIEHL24_14_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__16315\,
            in1 => \N__16834\,
            in2 => \N__16370\,
            in3 => \N__16792\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16524\,
            in2 => \_gnd_net_\,
            in3 => \N__16548\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_8_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16425\,
            in1 => \N__16449\,
            in2 => \N__16399\,
            in3 => \N__16467\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7KIH1_10_LC_8_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__16468\,
            in1 => \N__16293\,
            in2 => \N__18892\,
            in3 => \N__16493\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNISORB1_11_LC_8_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16549\,
            in1 => \N__16426\,
            in2 => \N__16531\,
            in3 => \N__16450\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2ALD3_14_LC_8_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__16331\,
            in1 => \N__16833\,
            in2 => \N__16325\,
            in3 => \N__16797\,
            lcout => \delay_measurement_inst.delay_hc_timer.un2_elapsed_time_hclto30_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_8_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16690\,
            in1 => \N__16747\,
            in2 => \N__16666\,
            in3 => \N__16717\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc_reg3lto19_3_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_8_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18847\,
            in2 => \N__18805\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_8_26_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_8_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18826\,
            in2 => \N__18781\,
            in3 => \N__16250\,
            lcout => \delay_measurement_inst.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_8_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18756\,
            in2 => \N__18806\,
            in3 => \N__16580\,
            lcout => \delay_measurement_inst.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_8_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19314\,
            in2 => \N__18782\,
            in3 => \N__16556\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_8_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18757\,
            in2 => \N__19297\,
            in3 => \N__16535\,
            lcout => \delay_measurement_inst.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_8_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19315\,
            in2 => \N__19273\,
            in3 => \N__16511\,
            lcout => \delay_measurement_inst.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_8_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19250\,
            in2 => \N__19298\,
            in3 => \N__16475\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_8_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19226\,
            in2 => \N__19274\,
            in3 => \N__16454\,
            lcout => \delay_measurement_inst.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__21973\,
            ce => \N__18868\,
            sr => \N__22295\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_8_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19249\,
            in2 => \N__19201\,
            in3 => \N__16430\,
            lcout => \delay_measurement_inst.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_8_27_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_8_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19225\,
            in2 => \N__19177\,
            in3 => \N__16403\,
            lcout => \delay_measurement_inst.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_8_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19152\,
            in2 => \N__19202\,
            in3 => \N__16373\,
            lcout => \delay_measurement_inst.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_8_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19134\,
            in2 => \N__19178\,
            in3 => \N__16802\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_8_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19153\,
            in2 => \N__19495\,
            in3 => \N__16754\,
            lcout => \delay_measurement_inst.delay_hc_reg3lto15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_8_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19135\,
            in2 => \N__19471\,
            in3 => \N__16724\,
            lcout => \delay_measurement_inst.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_8_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19448\,
            in2 => \N__19496\,
            in3 => \N__16697\,
            lcout => \delay_measurement_inst.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_8_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19424\,
            in2 => \N__19472\,
            in3 => \N__16670\,
            lcout => \delay_measurement_inst.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__21971\,
            ce => \N__18867\,
            sr => \N__22299\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_8_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19447\,
            in2 => \N__19399\,
            in3 => \N__16640\,
            lcout => \delay_measurement_inst.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_8_28_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_8_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19423\,
            in2 => \N__19375\,
            in3 => \N__16622\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_8_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19350\,
            in2 => \N__19400\,
            in3 => \N__16610\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_8_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19332\,
            in2 => \N__19376\,
            in3 => \N__16907\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_8_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19351\,
            in2 => \N__19684\,
            in3 => \N__16898\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_8_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19333\,
            in2 => \N__19660\,
            in3 => \N__16889\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_8_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19637\,
            in2 => \N__19685\,
            in3 => \N__16880\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_8_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19613\,
            in2 => \N__19661\,
            in3 => \N__16868\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__21967\,
            ce => \N__18866\,
            sr => \N__22302\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_8_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19636\,
            in2 => \N__19588\,
            in3 => \N__16859\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_8_29_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__21963\,
            ce => \N__18865\,
            sr => \N__22304\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_8_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19612\,
            in2 => \N__19564\,
            in3 => \N__16850\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__21963\,
            ce => \N__18865\,
            sr => \N__22304\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_8_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19540\,
            in2 => \N__19589\,
            in3 => \N__16841\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__21963\,
            ce => \N__18865\,
            sr => \N__22304\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_8_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19522\,
            in2 => \N__19565\,
            in3 => \N__17102\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__21963\,
            ce => \N__18865\,
            sr => \N__22304\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_8_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17099\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21963\,
            ce => \N__18865\,
            sr => \N__22304\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17072\,
            in2 => \N__17051\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17036\,
            in2 => \_gnd_net_\,
            in3 => \N__17018\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17015\,
            in2 => \N__17003\,
            in3 => \N__16985\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16982\,
            in2 => \_gnd_net_\,
            in3 => \N__16964\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16961\,
            in2 => \_gnd_net_\,
            in3 => \N__16943\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16940\,
            in2 => \_gnd_net_\,
            in3 => \N__16922\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17291\,
            in2 => \_gnd_net_\,
            in3 => \N__17273\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17270\,
            in2 => \_gnd_net_\,
            in3 => \N__17252\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17249\,
            in2 => \_gnd_net_\,
            in3 => \N__17231\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17228\,
            in2 => \_gnd_net_\,
            in3 => \N__17207\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17204\,
            in2 => \_gnd_net_\,
            in3 => \N__17186\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17179\,
            in2 => \_gnd_net_\,
            in3 => \N__17159\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17156\,
            in2 => \_gnd_net_\,
            in3 => \N__17135\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17132\,
            in2 => \_gnd_net_\,
            in3 => \N__17114\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17669\,
            in2 => \_gnd_net_\,
            in3 => \N__17648\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17645\,
            in2 => \_gnd_net_\,
            in3 => \N__17627\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17624\,
            in2 => \_gnd_net_\,
            in3 => \N__17606\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17603\,
            in2 => \_gnd_net_\,
            in3 => \N__17585\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17582\,
            in2 => \_gnd_net_\,
            in3 => \N__17570\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.stoper_state_0_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__17507\,
            in1 => \N__17398\,
            in2 => \N__20812\,
            in3 => \N__19714\,
            lcout => \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22005\,
            ce => \N__21342\,
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18422\,
            in2 => \N__17327\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_17_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17312\,
            in2 => \_gnd_net_\,
            in3 => \N__17294\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17867\,
            in2 => \N__17855\,
            in3 => \N__17831\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17828\,
            in2 => \_gnd_net_\,
            in3 => \N__17810\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17807\,
            in2 => \_gnd_net_\,
            in3 => \N__17789\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17786\,
            in2 => \_gnd_net_\,
            in3 => \N__17768\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17765\,
            in2 => \_gnd_net_\,
            in3 => \N__17747\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17744\,
            in2 => \_gnd_net_\,
            in3 => \N__17714\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17711\,
            in2 => \_gnd_net_\,
            in3 => \N__17693\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_18_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17690\,
            in2 => \_gnd_net_\,
            in3 => \N__17672\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18032\,
            in2 => \_gnd_net_\,
            in3 => \N__18014\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18011\,
            in2 => \_gnd_net_\,
            in3 => \N__17993\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17990\,
            in2 => \_gnd_net_\,
            in3 => \N__17972\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17969\,
            in2 => \_gnd_net_\,
            in3 => \N__17951\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17948\,
            in2 => \_gnd_net_\,
            in3 => \N__17930\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17926\,
            in2 => \_gnd_net_\,
            in3 => \N__17906\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17903\,
            in2 => \_gnd_net_\,
            in3 => \N__17882\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17879\,
            in2 => \_gnd_net_\,
            in3 => \N__18524\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18521\,
            in2 => \_gnd_net_\,
            in3 => \N__18509\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__18215\,
            in1 => \N__20523\,
            in2 => \_gnd_net_\,
            in3 => \N__18347\,
            lcout => \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18446\,
            in1 => \N__18418\,
            in2 => \_gnd_net_\,
            in3 => \N__18398\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20285\,
            in2 => \_gnd_net_\,
            in3 => \N__20365\,
            lcout => \phase_controller_slave.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20545\,
            in1 => \N__18321\,
            in2 => \_gnd_net_\,
            in3 => \N__18216\,
            lcout => \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_hc_RNO_0_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21222\,
            in2 => \_gnd_net_\,
            in3 => \N__21203\,
            lcout => \phase_controller_slave.N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.S1_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20288\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21984\,
            ce => 'H',
            sr => \N__22265\
        );

    \phase_controller_slave.stoper_hc.time_passed_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010101100"
        )
    port map (
            in0 => \N__21205\,
            in1 => \N__18110\,
            in2 => \N__18077\,
            in3 => \N__18062\,
            lcout => \phase_controller_slave.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21984\,
            ce => 'H',
            sr => \N__22265\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_14_5_LC_9_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18622\,
            in1 => \N__18634\,
            in2 => \N__18674\,
            in3 => \N__18544\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un2_startlto30_14_4_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18646\,
            in1 => \N__18658\,
            in2 => \N__18929\,
            in3 => \N__18556\,
            lcout => \phase_controller_inst1.stoper_hc.un2_startlto30_14Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_reg_30_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__18609\,
            in1 => \_gnd_net_\,
            in2 => \N__19117\,
            in3 => \N__18673\,
            lcout => measured_delay_hc_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_24_LC_9_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18659\,
            in1 => \N__19073\,
            in2 => \_gnd_net_\,
            in3 => \N__18985\,
            lcout => measured_delay_hc_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_25_LC_9_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__18986\,
            in1 => \_gnd_net_\,
            in2 => \N__19114\,
            in3 => \N__18647\,
            lcout => measured_delay_hc_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_28_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18635\,
            in1 => \N__19081\,
            in2 => \_gnd_net_\,
            in3 => \N__18989\,
            lcout => measured_delay_hc_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_29_LC_9_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__18608\,
            in1 => \_gnd_net_\,
            in2 => \N__19116\,
            in3 => \N__18623\,
            lcout => measured_delay_hc_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_23_LC_9_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__18557\,
            in1 => \N__18607\,
            in2 => \_gnd_net_\,
            in3 => \N__19072\,
            lcout => measured_delay_hc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_27_LC_9_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__18988\,
            in1 => \_gnd_net_\,
            in2 => \N__19115\,
            in3 => \N__18545\,
            lcout => measured_delay_hc_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_reg_26_LC_9_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18928\,
            in1 => \N__19077\,
            in2 => \_gnd_net_\,
            in3 => \N__18987\,
            lcout => measured_delay_hc_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21976\,
            ce => 'H',
            sr => \N__22283\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_9_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18848\,
            lcout => \delay_measurement_inst.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21974\,
            ce => \N__18869\,
            sr => \N__22287\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_9_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18827\,
            lcout => \delay_measurement_inst.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21974\,
            ce => \N__18869\,
            sr => \N__22287\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21034\,
            in1 => \N__18846\,
            in2 => \_gnd_net_\,
            in3 => \N__18830\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_26_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21059\,
            in1 => \N__18825\,
            in2 => \_gnd_net_\,
            in3 => \N__18809\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21035\,
            in1 => \N__18804\,
            in2 => \_gnd_net_\,
            in3 => \N__18785\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21060\,
            in1 => \N__18780\,
            in2 => \_gnd_net_\,
            in3 => \N__18761\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21036\,
            in1 => \N__18758\,
            in2 => \_gnd_net_\,
            in3 => \N__18743\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21061\,
            in1 => \N__19316\,
            in2 => \_gnd_net_\,
            in3 => \N__19301\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21037\,
            in1 => \N__19296\,
            in2 => \_gnd_net_\,
            in3 => \N__19277\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21062\,
            in1 => \N__19272\,
            in2 => \_gnd_net_\,
            in3 => \N__19253\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__21972\,
            ce => \N__21596\,
            sr => \N__22292\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21041\,
            in1 => \N__19248\,
            in2 => \_gnd_net_\,
            in3 => \N__19229\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_27_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21045\,
            in1 => \N__19224\,
            in2 => \_gnd_net_\,
            in3 => \N__19205\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21038\,
            in1 => \N__19200\,
            in2 => \_gnd_net_\,
            in3 => \N__19181\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21042\,
            in1 => \N__19176\,
            in2 => \_gnd_net_\,
            in3 => \N__19157\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21039\,
            in1 => \N__19154\,
            in2 => \_gnd_net_\,
            in3 => \N__19139\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21043\,
            in1 => \N__19136\,
            in2 => \_gnd_net_\,
            in3 => \N__19121\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21040\,
            in1 => \N__19494\,
            in2 => \_gnd_net_\,
            in3 => \N__19475\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21044\,
            in1 => \N__19470\,
            in2 => \_gnd_net_\,
            in3 => \N__19451\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__21968\,
            ce => \N__21606\,
            sr => \N__22296\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21072\,
            in1 => \N__19446\,
            in2 => \_gnd_net_\,
            in3 => \N__19427\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_9_28_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21055\,
            in1 => \N__19422\,
            in2 => \_gnd_net_\,
            in3 => \N__19403\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21073\,
            in1 => \N__19398\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21056\,
            in1 => \N__19374\,
            in2 => \_gnd_net_\,
            in3 => \N__19355\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21074\,
            in1 => \N__19352\,
            in2 => \_gnd_net_\,
            in3 => \N__19337\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21057\,
            in1 => \N__19334\,
            in2 => \_gnd_net_\,
            in3 => \N__19319\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21075\,
            in1 => \N__19683\,
            in2 => \_gnd_net_\,
            in3 => \N__19664\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21058\,
            in1 => \N__19659\,
            in2 => \_gnd_net_\,
            in3 => \N__19640\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__21964\,
            ce => \N__21607\,
            sr => \N__22300\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21063\,
            in1 => \N__19635\,
            in2 => \_gnd_net_\,
            in3 => \N__19616\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_9_29_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__21961\,
            ce => \N__21608\,
            sr => \N__22303\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21076\,
            in1 => \N__19611\,
            in2 => \_gnd_net_\,
            in3 => \N__19592\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__21961\,
            ce => \N__21608\,
            sr => \N__22303\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21064\,
            in1 => \N__19587\,
            in2 => \_gnd_net_\,
            in3 => \N__19568\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__21961\,
            ce => \N__21608\,
            sr => \N__22303\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21077\,
            in1 => \N__19563\,
            in2 => \_gnd_net_\,
            in3 => \N__19544\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__21961\,
            ce => \N__21608\,
            sr => \N__22303\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__21065\,
            in1 => \N__19541\,
            in2 => \_gnd_net_\,
            in3 => \N__19529\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__21961\,
            ce => \N__21608\,
            sr => \N__22303\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__19523\,
            in1 => \N__21066\,
            in2 => \_gnd_net_\,
            in3 => \N__19526\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21961\,
            ce => \N__21608\,
            sr => \N__22303\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21513\,
            in2 => \_gnd_net_\,
            in3 => \N__21479\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_138_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D1_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \il_max_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22017\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MAX_D2_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20168\,
            lcout => \il_max_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22011\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20162\,
            lcout => \il_min_comp1_D1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH1_MIN_D2_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20144\,
            lcout => \il_min_comp1_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22007\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20138\,
            in2 => \_gnd_net_\,
            in3 => \N__20033\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21999\,
            ce => \N__19945\,
            sr => \N__22232\
        );

    \phase_controller_inst1.state_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__21181\,
            in1 => \N__20249\,
            in2 => \N__20267\,
            in3 => \N__20209\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21994\,
            ce => 'H',
            sr => \N__22235\
        );

    \phase_controller_slave.start_timer_tr_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__19788\,
            in1 => \N__20237\,
            in2 => \N__20344\,
            in3 => \N__20216\,
            lcout => \phase_controller_slave.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21994\,
            ce => 'H',
            sr => \N__22235\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010100010111000"
        )
    port map (
            in0 => \N__20266\,
            in1 => \N__19751\,
            in2 => \N__19742\,
            in3 => \N__19718\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21994\,
            ce => 'H',
            sr => \N__22235\
        );

    \phase_controller_inst1.state_RNI7NN7_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20262\,
            in2 => \_gnd_net_\,
            in3 => \N__20248\,
            lcout => \phase_controller_inst1.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNIR0JF_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21170\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20208\,
            lcout => \phase_controller_inst1.T01_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_RNO_1_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21125\,
            in2 => \_gnd_net_\,
            in3 => \N__21240\,
            lcout => \phase_controller_slave.start_timer_tr_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_PH2_MIN_D2_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20231\,
            lcout => \il_min_comp2_D2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21991\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_1_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21548\,
            in2 => \_gnd_net_\,
            in3 => \N__20679\,
            lcout => \phase_controller_inst1.start_timer_hc_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.start_timer_tr_RNO_0_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20496\,
            in2 => \_gnd_net_\,
            in3 => \N__20463\,
            lcout => \phase_controller_slave.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__20438\,
            in1 => \N__20417\,
            in2 => \N__21180\,
            in3 => \N__20210\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_slave.state_0_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__21248\,
            in1 => \N__20497\,
            in2 => \N__21131\,
            in3 => \N__20464\,
            lcout => \phase_controller_slave.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_inst1.state_2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__20681\,
            in1 => \N__20436\,
            in2 => \N__21556\,
            in3 => \N__20416\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_inst1.T01_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__20437\,
            in1 => \N__20450\,
            in2 => \N__21644\,
            in3 => \N__20854\,
            lcout => shift_flag_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_inst1.start_timer_tr_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__20855\,
            in1 => \N__21643\,
            in2 => \N__20778\,
            in3 => \N__20689\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_inst1.state_3_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__20690\,
            in1 => \N__21552\,
            in2 => \N__21617\,
            in3 => \N__20680\,
            lcout => \phase_controller_inst1.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_inst1.start_timer_hc_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__20663\,
            in1 => \N__21642\,
            in2 => \N__20594\,
            in3 => \N__20381\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_slave.state_4_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__20299\,
            in1 => \N__20498\,
            in2 => \N__20333\,
            in3 => \N__20465\,
            lcout => \phase_controller_slave.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21987\,
            ce => 'H',
            sr => \N__22240\
        );

    \phase_controller_slave.un1_start_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21709\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20449\,
            lcout => \phase_controller_slave.un1_startZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_hc_RNO_0_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20435\,
            in2 => \_gnd_net_\,
            in3 => \N__20410\,
            lcout => \phase_controller_inst1.N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_slave.state_2_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__20375\,
            in1 => \N__20287\,
            in2 => \N__21227\,
            in3 => \N__21204\,
            lcout => \phase_controller_slave.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21981\,
            ce => 'H',
            sr => \N__22247\
        );

    \phase_controller_slave.state_3_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001000000010"
        )
    port map (
            in0 => \N__20286\,
            in1 => \N__20374\,
            in2 => \N__20343\,
            in3 => \N__20300\,
            lcout => \phase_controller_slave.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21981\,
            ce => 'H',
            sr => \N__22247\
        );

    \phase_controller_slave.state_1_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__21247\,
            in1 => \N__21226\,
            in2 => \N__21126\,
            in3 => \N__21206\,
            lcout => \phase_controller_slave.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21978\,
            ce => 'H',
            sr => \N__22252\
        );

    \phase_controller_inst1.S2_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21182\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21977\,
            ce => 'H',
            sr => \N__22259\
        );

    \phase_controller_slave.S2_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21130\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21969\,
            ce => 'H',
            sr => \N__22277\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21761\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__21515\,
            in1 => \N__21497\,
            in2 => \_gnd_net_\,
            in3 => \N__21484\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22012\,
            ce => 'H',
            sr => \N__22231\
        );

    \delay_measurement_inst.stop_timer_tr_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21394\,
            in1 => \N__21419\,
            in2 => \_gnd_net_\,
            in3 => \N__21374\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22012\,
            ce => 'H',
            sr => \N__22231\
        );

    \delay_measurement_inst.start_timer_tr_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21418\,
            in1 => \N__21373\,
            in2 => \_gnd_net_\,
            in3 => \N__21393\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22012\,
            ce => 'H',
            sr => \N__22231\
        );

    \delay_measurement_inst.prev_tr_sig_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21420\,
            lcout => \delay_measurement_inst.prev_tr_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22012\,
            ce => 'H',
            sr => \N__22231\
        );

    \delay_measurement_inst.tr_state_RNIFBI31_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__21371\,
            in1 => \N__21392\,
            in2 => \N__21422\,
            in3 => \N__20951\,
            lcout => \delay_measurement_inst.un1_tr_state_1_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_4_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21707\,
            in2 => \_gnd_net_\,
            in3 => \N__21638\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21988\,
            ce => 'H',
            sr => \N__22236\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21637\,
            lcout => \phase_controller_inst1.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_11_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__22414\,
            in1 => \N__21785\,
            in2 => \_gnd_net_\,
            in3 => \N__21759\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_137_i_g\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S1_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21563\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21959\,
            ce => 'H',
            sr => \N__22288\
        );

    \SB_DFF_inst_DELAY_TR2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21428\,
            lcout => delay_tr_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__21514\,
            in1 => \N__21496\,
            in2 => \_gnd_net_\,
            in3 => \N__21480\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_139_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_TR1_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21446\,
            lcout => delay_tr_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22006\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.tr_state_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__21372\,
            in2 => \_gnd_net_\,
            in3 => \N__21395\,
            lcout => \delay_measurement_inst.tr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21998\,
            ce => \N__21349\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.hc_state_0_LC_12_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__22377\,
            in1 => \N__22359\,
            in2 => \_gnd_net_\,
            in3 => \N__22071\,
            lcout => \delay_measurement_inst.hc_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21965\,
            ce => \N__21338\,
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.start_timer_hc_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__22379\,
            in1 => \N__22360\,
            in2 => \_gnd_net_\,
            in3 => \N__22076\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21962\,
            ce => 'H',
            sr => \N__22269\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_12_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__22415\,
            in1 => \N__21781\,
            in2 => \_gnd_net_\,
            in3 => \N__21760\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21960\,
            ce => 'H',
            sr => \N__22274\
        );

    \SB_DFF_inst_DELAY_HC1_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => delay_hc_d1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SB_DFF_inst_DELAY_HC2_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22388\,
            lcout => delay_hc_d2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.prev_hc_sig_LC_13_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22075\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.prev_hc_sigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21970\,
            ce => 'H',
            sr => \N__22253\
        );

    \delay_measurement_inst.stop_timer_hc_LC_13_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__22378\,
            in1 => \N__22361\,
            in2 => \N__22343\,
            in3 => \N__22070\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21777\,
            in2 => \_gnd_net_\,
            in3 => \N__21755\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_136_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
