// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 15 2025 13:11:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    start_stop,
    s2_phy,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    input start_stop;
    output s2_phy;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__47202;
    wire N__47201;
    wire N__47200;
    wire N__47191;
    wire N__47190;
    wire N__47189;
    wire N__47182;
    wire N__47181;
    wire N__47180;
    wire N__47173;
    wire N__47172;
    wire N__47171;
    wire N__47164;
    wire N__47163;
    wire N__47162;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47146;
    wire N__47145;
    wire N__47144;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47128;
    wire N__47127;
    wire N__47126;
    wire N__47119;
    wire N__47118;
    wire N__47117;
    wire N__47110;
    wire N__47109;
    wire N__47108;
    wire N__47101;
    wire N__47100;
    wire N__47099;
    wire N__47092;
    wire N__47091;
    wire N__47090;
    wire N__47073;
    wire N__47070;
    wire N__47069;
    wire N__47066;
    wire N__47063;
    wire N__47062;
    wire N__47061;
    wire N__47060;
    wire N__47059;
    wire N__47056;
    wire N__47053;
    wire N__47044;
    wire N__47041;
    wire N__47038;
    wire N__47035;
    wire N__47028;
    wire N__47025;
    wire N__47022;
    wire N__47021;
    wire N__47020;
    wire N__47017;
    wire N__47014;
    wire N__47011;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46984;
    wire N__46983;
    wire N__46982;
    wire N__46979;
    wire N__46976;
    wire N__46973;
    wire N__46970;
    wire N__46967;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46943;
    wire N__46942;
    wire N__46941;
    wire N__46940;
    wire N__46939;
    wire N__46938;
    wire N__46937;
    wire N__46936;
    wire N__46935;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46912;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46896;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46890;
    wire N__46873;
    wire N__46868;
    wire N__46853;
    wire N__46850;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46837;
    wire N__46836;
    wire N__46835;
    wire N__46834;
    wire N__46833;
    wire N__46832;
    wire N__46831;
    wire N__46830;
    wire N__46829;
    wire N__46828;
    wire N__46825;
    wire N__46822;
    wire N__46815;
    wire N__46808;
    wire N__46805;
    wire N__46792;
    wire N__46791;
    wire N__46784;
    wire N__46781;
    wire N__46776;
    wire N__46769;
    wire N__46766;
    wire N__46755;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46747;
    wire N__46746;
    wire N__46743;
    wire N__46740;
    wire N__46735;
    wire N__46734;
    wire N__46733;
    wire N__46732;
    wire N__46731;
    wire N__46730;
    wire N__46729;
    wire N__46726;
    wire N__46721;
    wire N__46718;
    wire N__46717;
    wire N__46716;
    wire N__46715;
    wire N__46714;
    wire N__46713;
    wire N__46712;
    wire N__46703;
    wire N__46702;
    wire N__46701;
    wire N__46698;
    wire N__46693;
    wire N__46686;
    wire N__46681;
    wire N__46678;
    wire N__46675;
    wire N__46672;
    wire N__46667;
    wire N__46664;
    wire N__46647;
    wire N__46644;
    wire N__46643;
    wire N__46642;
    wire N__46641;
    wire N__46638;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46607;
    wire N__46602;
    wire N__46593;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46578;
    wire N__46577;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46565;
    wire N__46562;
    wire N__46561;
    wire N__46558;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46535;
    wire N__46528;
    wire N__46523;
    wire N__46520;
    wire N__46515;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46505;
    wire N__46500;
    wire N__46499;
    wire N__46498;
    wire N__46497;
    wire N__46496;
    wire N__46495;
    wire N__46494;
    wire N__46493;
    wire N__46492;
    wire N__46491;
    wire N__46488;
    wire N__46485;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46481;
    wire N__46478;
    wire N__46475;
    wire N__46474;
    wire N__46473;
    wire N__46470;
    wire N__46469;
    wire N__46466;
    wire N__46465;
    wire N__46462;
    wire N__46461;
    wire N__46460;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46452;
    wire N__46451;
    wire N__46450;
    wire N__46449;
    wire N__46440;
    wire N__46439;
    wire N__46434;
    wire N__46423;
    wire N__46414;
    wire N__46409;
    wire N__46406;
    wire N__46395;
    wire N__46392;
    wire N__46389;
    wire N__46388;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46380;
    wire N__46379;
    wire N__46378;
    wire N__46375;
    wire N__46370;
    wire N__46367;
    wire N__46362;
    wire N__46353;
    wire N__46352;
    wire N__46347;
    wire N__46340;
    wire N__46335;
    wire N__46328;
    wire N__46325;
    wire N__46320;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46304;
    wire N__46301;
    wire N__46298;
    wire N__46293;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46281;
    wire N__46280;
    wire N__46279;
    wire N__46278;
    wire N__46277;
    wire N__46276;
    wire N__46275;
    wire N__46274;
    wire N__46273;
    wire N__46272;
    wire N__46271;
    wire N__46270;
    wire N__46269;
    wire N__46268;
    wire N__46267;
    wire N__46266;
    wire N__46265;
    wire N__46256;
    wire N__46255;
    wire N__46254;
    wire N__46253;
    wire N__46252;
    wire N__46251;
    wire N__46250;
    wire N__46249;
    wire N__46248;
    wire N__46243;
    wire N__46232;
    wire N__46223;
    wire N__46222;
    wire N__46221;
    wire N__46220;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46193;
    wire N__46190;
    wire N__46185;
    wire N__46178;
    wire N__46177;
    wire N__46176;
    wire N__46175;
    wire N__46174;
    wire N__46171;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46153;
    wire N__46144;
    wire N__46131;
    wire N__46130;
    wire N__46129;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46112;
    wire N__46109;
    wire N__46106;
    wire N__46103;
    wire N__46100;
    wire N__46097;
    wire N__46094;
    wire N__46091;
    wire N__46086;
    wire N__46077;
    wire N__46076;
    wire N__46075;
    wire N__46074;
    wire N__46073;
    wire N__46072;
    wire N__46071;
    wire N__46070;
    wire N__46069;
    wire N__46068;
    wire N__46067;
    wire N__46066;
    wire N__46065;
    wire N__46064;
    wire N__46063;
    wire N__46062;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46058;
    wire N__46057;
    wire N__46056;
    wire N__46055;
    wire N__46054;
    wire N__46053;
    wire N__46052;
    wire N__46051;
    wire N__46050;
    wire N__46049;
    wire N__46048;
    wire N__46047;
    wire N__46046;
    wire N__46045;
    wire N__46044;
    wire N__46043;
    wire N__46042;
    wire N__46041;
    wire N__46040;
    wire N__46039;
    wire N__46038;
    wire N__46037;
    wire N__46036;
    wire N__46035;
    wire N__46034;
    wire N__46033;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46028;
    wire N__46027;
    wire N__46026;
    wire N__46025;
    wire N__46024;
    wire N__46023;
    wire N__46022;
    wire N__46021;
    wire N__46020;
    wire N__46019;
    wire N__46018;
    wire N__46017;
    wire N__46016;
    wire N__46015;
    wire N__46014;
    wire N__46013;
    wire N__46012;
    wire N__46011;
    wire N__46010;
    wire N__46009;
    wire N__46008;
    wire N__46007;
    wire N__46006;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__46001;
    wire N__46000;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45990;
    wire N__45989;
    wire N__45988;
    wire N__45987;
    wire N__45986;
    wire N__45985;
    wire N__45984;
    wire N__45983;
    wire N__45982;
    wire N__45981;
    wire N__45980;
    wire N__45979;
    wire N__45978;
    wire N__45977;
    wire N__45976;
    wire N__45975;
    wire N__45974;
    wire N__45973;
    wire N__45972;
    wire N__45971;
    wire N__45970;
    wire N__45969;
    wire N__45968;
    wire N__45967;
    wire N__45966;
    wire N__45965;
    wire N__45964;
    wire N__45963;
    wire N__45962;
    wire N__45961;
    wire N__45960;
    wire N__45959;
    wire N__45958;
    wire N__45957;
    wire N__45956;
    wire N__45955;
    wire N__45954;
    wire N__45953;
    wire N__45952;
    wire N__45951;
    wire N__45950;
    wire N__45949;
    wire N__45948;
    wire N__45947;
    wire N__45946;
    wire N__45945;
    wire N__45944;
    wire N__45943;
    wire N__45942;
    wire N__45941;
    wire N__45940;
    wire N__45939;
    wire N__45938;
    wire N__45937;
    wire N__45936;
    wire N__45935;
    wire N__45934;
    wire N__45933;
    wire N__45932;
    wire N__45931;
    wire N__45930;
    wire N__45929;
    wire N__45928;
    wire N__45627;
    wire N__45624;
    wire N__45623;
    wire N__45622;
    wire N__45621;
    wire N__45620;
    wire N__45619;
    wire N__45618;
    wire N__45615;
    wire N__45612;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45581;
    wire N__45580;
    wire N__45579;
    wire N__45578;
    wire N__45577;
    wire N__45576;
    wire N__45575;
    wire N__45574;
    wire N__45573;
    wire N__45572;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45566;
    wire N__45565;
    wire N__45564;
    wire N__45563;
    wire N__45562;
    wire N__45561;
    wire N__45560;
    wire N__45559;
    wire N__45558;
    wire N__45557;
    wire N__45556;
    wire N__45555;
    wire N__45554;
    wire N__45553;
    wire N__45552;
    wire N__45551;
    wire N__45550;
    wire N__45549;
    wire N__45548;
    wire N__45547;
    wire N__45546;
    wire N__45545;
    wire N__45544;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45540;
    wire N__45539;
    wire N__45536;
    wire N__45535;
    wire N__45534;
    wire N__45533;
    wire N__45532;
    wire N__45531;
    wire N__45530;
    wire N__45529;
    wire N__45528;
    wire N__45527;
    wire N__45526;
    wire N__45525;
    wire N__45524;
    wire N__45523;
    wire N__45522;
    wire N__45521;
    wire N__45520;
    wire N__45519;
    wire N__45518;
    wire N__45517;
    wire N__45516;
    wire N__45515;
    wire N__45514;
    wire N__45513;
    wire N__45512;
    wire N__45511;
    wire N__45510;
    wire N__45509;
    wire N__45508;
    wire N__45507;
    wire N__45506;
    wire N__45505;
    wire N__45504;
    wire N__45503;
    wire N__45502;
    wire N__45501;
    wire N__45500;
    wire N__45499;
    wire N__45498;
    wire N__45497;
    wire N__45496;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45492;
    wire N__45491;
    wire N__45490;
    wire N__45489;
    wire N__45488;
    wire N__45487;
    wire N__45486;
    wire N__45485;
    wire N__45484;
    wire N__45483;
    wire N__45482;
    wire N__45481;
    wire N__45480;
    wire N__45479;
    wire N__45478;
    wire N__45477;
    wire N__45476;
    wire N__45475;
    wire N__45474;
    wire N__45473;
    wire N__45470;
    wire N__45469;
    wire N__45468;
    wire N__45467;
    wire N__45466;
    wire N__45465;
    wire N__45462;
    wire N__45461;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45449;
    wire N__45448;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45440;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45149;
    wire N__45146;
    wire N__45143;
    wire N__45140;
    wire N__45137;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45068;
    wire N__45065;
    wire N__45062;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45023;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45009;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44973;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44957;
    wire N__44954;
    wire N__44951;
    wire N__44948;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44927;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44900;
    wire N__44897;
    wire N__44894;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44879;
    wire N__44876;
    wire N__44873;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44846;
    wire N__44843;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44814;
    wire N__44813;
    wire N__44810;
    wire N__44807;
    wire N__44804;
    wire N__44801;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44774;
    wire N__44771;
    wire N__44768;
    wire N__44765;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44708;
    wire N__44705;
    wire N__44702;
    wire N__44699;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44667;
    wire N__44666;
    wire N__44665;
    wire N__44664;
    wire N__44663;
    wire N__44662;
    wire N__44657;
    wire N__44654;
    wire N__44653;
    wire N__44650;
    wire N__44649;
    wire N__44648;
    wire N__44647;
    wire N__44646;
    wire N__44645;
    wire N__44644;
    wire N__44643;
    wire N__44642;
    wire N__44641;
    wire N__44640;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44632;
    wire N__44631;
    wire N__44628;
    wire N__44623;
    wire N__44606;
    wire N__44603;
    wire N__44600;
    wire N__44597;
    wire N__44586;
    wire N__44585;
    wire N__44584;
    wire N__44579;
    wire N__44576;
    wire N__44569;
    wire N__44566;
    wire N__44561;
    wire N__44560;
    wire N__44559;
    wire N__44554;
    wire N__44547;
    wire N__44544;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44511;
    wire N__44510;
    wire N__44509;
    wire N__44508;
    wire N__44507;
    wire N__44506;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44490;
    wire N__44489;
    wire N__44486;
    wire N__44483;
    wire N__44482;
    wire N__44481;
    wire N__44478;
    wire N__44477;
    wire N__44476;
    wire N__44475;
    wire N__44474;
    wire N__44473;
    wire N__44472;
    wire N__44455;
    wire N__44446;
    wire N__44445;
    wire N__44444;
    wire N__44441;
    wire N__44434;
    wire N__44433;
    wire N__44430;
    wire N__44429;
    wire N__44428;
    wire N__44423;
    wire N__44418;
    wire N__44413;
    wire N__44410;
    wire N__44407;
    wire N__44404;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44380;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44357;
    wire N__44354;
    wire N__44353;
    wire N__44352;
    wire N__44351;
    wire N__44350;
    wire N__44349;
    wire N__44348;
    wire N__44347;
    wire N__44346;
    wire N__44345;
    wire N__44344;
    wire N__44343;
    wire N__44342;
    wire N__44341;
    wire N__44340;
    wire N__44339;
    wire N__44338;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44314;
    wire N__44303;
    wire N__44302;
    wire N__44301;
    wire N__44300;
    wire N__44299;
    wire N__44298;
    wire N__44295;
    wire N__44288;
    wire N__44283;
    wire N__44278;
    wire N__44275;
    wire N__44268;
    wire N__44263;
    wire N__44252;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44221;
    wire N__44218;
    wire N__44215;
    wire N__44212;
    wire N__44207;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44180;
    wire N__44177;
    wire N__44174;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44156;
    wire N__44153;
    wire N__44150;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43952;
    wire N__43949;
    wire N__43946;
    wire N__43945;
    wire N__43944;
    wire N__43941;
    wire N__43936;
    wire N__43933;
    wire N__43928;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43880;
    wire N__43877;
    wire N__43874;
    wire N__43871;
    wire N__43870;
    wire N__43867;
    wire N__43864;
    wire N__43861;
    wire N__43854;
    wire N__43851;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43841;
    wire N__43838;
    wire N__43833;
    wire N__43830;
    wire N__43829;
    wire N__43828;
    wire N__43827;
    wire N__43826;
    wire N__43825;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43805;
    wire N__43802;
    wire N__43801;
    wire N__43798;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43776;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43762;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43750;
    wire N__43747;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43731;
    wire N__43730;
    wire N__43729;
    wire N__43728;
    wire N__43723;
    wire N__43722;
    wire N__43721;
    wire N__43716;
    wire N__43713;
    wire N__43708;
    wire N__43707;
    wire N__43706;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43691;
    wire N__43688;
    wire N__43677;
    wire N__43676;
    wire N__43675;
    wire N__43674;
    wire N__43673;
    wire N__43672;
    wire N__43671;
    wire N__43670;
    wire N__43667;
    wire N__43666;
    wire N__43665;
    wire N__43662;
    wire N__43661;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43649;
    wire N__43648;
    wire N__43647;
    wire N__43636;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43615;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43590;
    wire N__43581;
    wire N__43578;
    wire N__43577;
    wire N__43576;
    wire N__43573;
    wire N__43568;
    wire N__43565;
    wire N__43562;
    wire N__43557;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43543;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43531;
    wire N__43524;
    wire N__43521;
    wire N__43520;
    wire N__43519;
    wire N__43516;
    wire N__43515;
    wire N__43512;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43480;
    wire N__43473;
    wire N__43472;
    wire N__43471;
    wire N__43470;
    wire N__43469;
    wire N__43468;
    wire N__43455;
    wire N__43454;
    wire N__43453;
    wire N__43452;
    wire N__43451;
    wire N__43450;
    wire N__43449;
    wire N__43448;
    wire N__43447;
    wire N__43446;
    wire N__43445;
    wire N__43444;
    wire N__43443;
    wire N__43442;
    wire N__43439;
    wire N__43430;
    wire N__43429;
    wire N__43428;
    wire N__43425;
    wire N__43412;
    wire N__43407;
    wire N__43402;
    wire N__43401;
    wire N__43398;
    wire N__43397;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43363;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43341;
    wire N__43340;
    wire N__43339;
    wire N__43338;
    wire N__43337;
    wire N__43336;
    wire N__43335;
    wire N__43334;
    wire N__43333;
    wire N__43332;
    wire N__43331;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43317;
    wire N__43316;
    wire N__43315;
    wire N__43312;
    wire N__43311;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43292;
    wire N__43291;
    wire N__43290;
    wire N__43287;
    wire N__43286;
    wire N__43285;
    wire N__43284;
    wire N__43283;
    wire N__43270;
    wire N__43265;
    wire N__43256;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43234;
    wire N__43231;
    wire N__43228;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43216;
    wire N__43211;
    wire N__43208;
    wire N__43205;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43187;
    wire N__43176;
    wire N__43173;
    wire N__43172;
    wire N__43169;
    wire N__43166;
    wire N__43165;
    wire N__43160;
    wire N__43157;
    wire N__43156;
    wire N__43155;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43133;
    wire N__43128;
    wire N__43127;
    wire N__43126;
    wire N__43125;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43117;
    wire N__43116;
    wire N__43115;
    wire N__43114;
    wire N__43111;
    wire N__43110;
    wire N__43109;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43101;
    wire N__43100;
    wire N__43099;
    wire N__43098;
    wire N__43093;
    wire N__43084;
    wire N__43083;
    wire N__43080;
    wire N__43073;
    wire N__43072;
    wire N__43071;
    wire N__43070;
    wire N__43069;
    wire N__43062;
    wire N__43055;
    wire N__43050;
    wire N__43047;
    wire N__43046;
    wire N__43043;
    wire N__43040;
    wire N__43035;
    wire N__43032;
    wire N__43031;
    wire N__43028;
    wire N__43023;
    wire N__43018;
    wire N__43015;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42996;
    wire N__42993;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42971;
    wire N__42960;
    wire N__42959;
    wire N__42958;
    wire N__42957;
    wire N__42956;
    wire N__42955;
    wire N__42954;
    wire N__42953;
    wire N__42952;
    wire N__42951;
    wire N__42950;
    wire N__42949;
    wire N__42948;
    wire N__42947;
    wire N__42944;
    wire N__42943;
    wire N__42940;
    wire N__42939;
    wire N__42938;
    wire N__42937;
    wire N__42936;
    wire N__42935;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42918;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42889;
    wire N__42872;
    wire N__42867;
    wire N__42864;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42849;
    wire N__42848;
    wire N__42839;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42814;
    wire N__42813;
    wire N__42812;
    wire N__42809;
    wire N__42808;
    wire N__42807;
    wire N__42806;
    wire N__42805;
    wire N__42798;
    wire N__42797;
    wire N__42794;
    wire N__42793;
    wire N__42792;
    wire N__42791;
    wire N__42790;
    wire N__42789;
    wire N__42788;
    wire N__42787;
    wire N__42786;
    wire N__42785;
    wire N__42782;
    wire N__42781;
    wire N__42780;
    wire N__42777;
    wire N__42776;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42753;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42725;
    wire N__42714;
    wire N__42711;
    wire N__42704;
    wire N__42701;
    wire N__42694;
    wire N__42681;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42673;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42659;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42641;
    wire N__42630;
    wire N__42629;
    wire N__42628;
    wire N__42627;
    wire N__42626;
    wire N__42625;
    wire N__42624;
    wire N__42623;
    wire N__42622;
    wire N__42621;
    wire N__42620;
    wire N__42619;
    wire N__42618;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42610;
    wire N__42609;
    wire N__42608;
    wire N__42607;
    wire N__42606;
    wire N__42605;
    wire N__42604;
    wire N__42603;
    wire N__42600;
    wire N__42585;
    wire N__42582;
    wire N__42581;
    wire N__42574;
    wire N__42569;
    wire N__42552;
    wire N__42549;
    wire N__42544;
    wire N__42541;
    wire N__42540;
    wire N__42535;
    wire N__42526;
    wire N__42523;
    wire N__42520;
    wire N__42517;
    wire N__42510;
    wire N__42509;
    wire N__42508;
    wire N__42507;
    wire N__42506;
    wire N__42503;
    wire N__42502;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42490;
    wire N__42487;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42463;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42437;
    wire N__42434;
    wire N__42423;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42401;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42372;
    wire N__42371;
    wire N__42368;
    wire N__42365;
    wire N__42362;
    wire N__42359;
    wire N__42358;
    wire N__42353;
    wire N__42350;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42335;
    wire N__42332;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42318;
    wire N__42317;
    wire N__42314;
    wire N__42311;
    wire N__42306;
    wire N__42305;
    wire N__42302;
    wire N__42299;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42278;
    wire N__42277;
    wire N__42276;
    wire N__42273;
    wire N__42266;
    wire N__42261;
    wire N__42260;
    wire N__42259;
    wire N__42258;
    wire N__42257;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42242;
    wire N__42239;
    wire N__42232;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42220;
    wire N__42213;
    wire N__42210;
    wire N__42207;
    wire N__42204;
    wire N__42201;
    wire N__42198;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42179;
    wire N__42176;
    wire N__42173;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42101;
    wire N__42098;
    wire N__42095;
    wire N__42090;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42078;
    wire N__42077;
    wire N__42076;
    wire N__42073;
    wire N__42070;
    wire N__42067;
    wire N__42066;
    wire N__42063;
    wire N__42058;
    wire N__42055;
    wire N__42050;
    wire N__42045;
    wire N__42044;
    wire N__42041;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42019;
    wire N__42014;
    wire N__42011;
    wire N__42006;
    wire N__42005;
    wire N__42002;
    wire N__41999;
    wire N__41998;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41954;
    wire N__41953;
    wire N__41950;
    wire N__41945;
    wire N__41940;
    wire N__41937;
    wire N__41936;
    wire N__41935;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41921;
    wire N__41918;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41885;
    wire N__41884;
    wire N__41881;
    wire N__41878;
    wire N__41875;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41863;
    wire N__41860;
    wire N__41859;
    wire N__41858;
    wire N__41855;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41836;
    wire N__41829;
    wire N__41828;
    wire N__41827;
    wire N__41824;
    wire N__41821;
    wire N__41818;
    wire N__41817;
    wire N__41816;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41797;
    wire N__41794;
    wire N__41791;
    wire N__41788;
    wire N__41781;
    wire N__41780;
    wire N__41779;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41771;
    wire N__41770;
    wire N__41769;
    wire N__41768;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41754;
    wire N__41753;
    wire N__41752;
    wire N__41751;
    wire N__41750;
    wire N__41749;
    wire N__41748;
    wire N__41747;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41737;
    wire N__41736;
    wire N__41735;
    wire N__41734;
    wire N__41733;
    wire N__41726;
    wire N__41723;
    wire N__41708;
    wire N__41699;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41681;
    wire N__41670;
    wire N__41669;
    wire N__41668;
    wire N__41665;
    wire N__41660;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41645;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41637;
    wire N__41634;
    wire N__41629;
    wire N__41626;
    wire N__41623;
    wire N__41622;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41598;
    wire N__41595;
    wire N__41594;
    wire N__41593;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41573;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41557;
    wire N__41554;
    wire N__41549;
    wire N__41546;
    wire N__41541;
    wire N__41540;
    wire N__41539;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41525;
    wire N__41524;
    wire N__41523;
    wire N__41522;
    wire N__41521;
    wire N__41518;
    wire N__41501;
    wire N__41500;
    wire N__41499;
    wire N__41498;
    wire N__41497;
    wire N__41496;
    wire N__41495;
    wire N__41494;
    wire N__41493;
    wire N__41492;
    wire N__41489;
    wire N__41486;
    wire N__41483;
    wire N__41480;
    wire N__41477;
    wire N__41476;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41465;
    wire N__41464;
    wire N__41463;
    wire N__41462;
    wire N__41461;
    wire N__41460;
    wire N__41459;
    wire N__41458;
    wire N__41457;
    wire N__41456;
    wire N__41455;
    wire N__41452;
    wire N__41447;
    wire N__41442;
    wire N__41439;
    wire N__41430;
    wire N__41417;
    wire N__41412;
    wire N__41399;
    wire N__41396;
    wire N__41391;
    wire N__41376;
    wire N__41375;
    wire N__41374;
    wire N__41373;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41294;
    wire N__41293;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41282;
    wire N__41279;
    wire N__41276;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41258;
    wire N__41253;
    wire N__41252;
    wire N__41249;
    wire N__41246;
    wire N__41241;
    wire N__41240;
    wire N__41239;
    wire N__41238;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41225;
    wire N__41224;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41208;
    wire N__41203;
    wire N__41196;
    wire N__41195;
    wire N__41192;
    wire N__41191;
    wire N__41188;
    wire N__41187;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41163;
    wire N__41160;
    wire N__41151;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41123;
    wire N__41120;
    wire N__41119;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41098;
    wire N__41097;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41079;
    wire N__41076;
    wire N__41075;
    wire N__41072;
    wire N__41071;
    wire N__41070;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41054;
    wire N__41051;
    wire N__41046;
    wire N__41041;
    wire N__41034;
    wire N__41031;
    wire N__41030;
    wire N__41029;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41004;
    wire N__41001;
    wire N__40992;
    wire N__40991;
    wire N__40990;
    wire N__40987;
    wire N__40984;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40971;
    wire N__40970;
    wire N__40967;
    wire N__40962;
    wire N__40957;
    wire N__40950;
    wire N__40947;
    wire N__40946;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40938;
    wire N__40937;
    wire N__40934;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40918;
    wire N__40915;
    wire N__40912;
    wire N__40907;
    wire N__40902;
    wire N__40899;
    wire N__40898;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40886;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40865;
    wire N__40862;
    wire N__40859;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40842;
    wire N__40839;
    wire N__40838;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40797;
    wire N__40794;
    wire N__40793;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40782;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40768;
    wire N__40761;
    wire N__40760;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40749;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40733;
    wire N__40730;
    wire N__40727;
    wire N__40724;
    wire N__40719;
    wire N__40716;
    wire N__40715;
    wire N__40712;
    wire N__40709;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40692;
    wire N__40691;
    wire N__40688;
    wire N__40685;
    wire N__40684;
    wire N__40679;
    wire N__40676;
    wire N__40673;
    wire N__40668;
    wire N__40665;
    wire N__40664;
    wire N__40661;
    wire N__40658;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40643;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40628;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40605;
    wire N__40602;
    wire N__40601;
    wire N__40598;
    wire N__40595;
    wire N__40594;
    wire N__40589;
    wire N__40586;
    wire N__40583;
    wire N__40578;
    wire N__40575;
    wire N__40574;
    wire N__40573;
    wire N__40568;
    wire N__40565;
    wire N__40562;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40541;
    wire N__40536;
    wire N__40533;
    wire N__40532;
    wire N__40531;
    wire N__40530;
    wire N__40529;
    wire N__40528;
    wire N__40527;
    wire N__40526;
    wire N__40525;
    wire N__40524;
    wire N__40523;
    wire N__40522;
    wire N__40513;
    wire N__40504;
    wire N__40495;
    wire N__40494;
    wire N__40493;
    wire N__40492;
    wire N__40491;
    wire N__40490;
    wire N__40489;
    wire N__40488;
    wire N__40487;
    wire N__40486;
    wire N__40485;
    wire N__40478;
    wire N__40473;
    wire N__40464;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40460;
    wire N__40459;
    wire N__40458;
    wire N__40457;
    wire N__40456;
    wire N__40447;
    wire N__40440;
    wire N__40431;
    wire N__40422;
    wire N__40417;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40400;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40386;
    wire N__40385;
    wire N__40382;
    wire N__40379;
    wire N__40378;
    wire N__40377;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40358;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40314;
    wire N__40313;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40299;
    wire N__40296;
    wire N__40295;
    wire N__40292;
    wire N__40289;
    wire N__40288;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40272;
    wire N__40269;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40259;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40232;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40217;
    wire N__40212;
    wire N__40209;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40201;
    wire N__40196;
    wire N__40193;
    wire N__40190;
    wire N__40185;
    wire N__40182;
    wire N__40181;
    wire N__40178;
    wire N__40175;
    wire N__40170;
    wire N__40169;
    wire N__40166;
    wire N__40163;
    wire N__40160;
    wire N__40155;
    wire N__40152;
    wire N__40151;
    wire N__40148;
    wire N__40145;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40130;
    wire N__40125;
    wire N__40122;
    wire N__40121;
    wire N__40120;
    wire N__40115;
    wire N__40112;
    wire N__40109;
    wire N__40104;
    wire N__40101;
    wire N__40100;
    wire N__40099;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40083;
    wire N__40080;
    wire N__40079;
    wire N__40078;
    wire N__40073;
    wire N__40070;
    wire N__40067;
    wire N__40062;
    wire N__40059;
    wire N__40058;
    wire N__40055;
    wire N__40052;
    wire N__40047;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40032;
    wire N__40029;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40007;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39995;
    wire N__39992;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39977;
    wire N__39974;
    wire N__39969;
    wire N__39966;
    wire N__39965;
    wire N__39962;
    wire N__39959;
    wire N__39958;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39942;
    wire N__39939;
    wire N__39938;
    wire N__39937;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39921;
    wire N__39918;
    wire N__39917;
    wire N__39912;
    wire N__39911;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39890;
    wire N__39887;
    wire N__39886;
    wire N__39883;
    wire N__39880;
    wire N__39877;
    wire N__39872;
    wire N__39867;
    wire N__39864;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39856;
    wire N__39851;
    wire N__39848;
    wire N__39847;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39781;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39769;
    wire N__39762;
    wire N__39759;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39751;
    wire N__39746;
    wire N__39743;
    wire N__39740;
    wire N__39735;
    wire N__39732;
    wire N__39731;
    wire N__39730;
    wire N__39725;
    wire N__39722;
    wire N__39719;
    wire N__39714;
    wire N__39711;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39703;
    wire N__39700;
    wire N__39697;
    wire N__39694;
    wire N__39689;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39677;
    wire N__39674;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39664;
    wire N__39659;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39647;
    wire N__39644;
    wire N__39641;
    wire N__39638;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39504;
    wire N__39503;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39479;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39465;
    wire N__39464;
    wire N__39461;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39441;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39429;
    wire N__39426;
    wire N__39425;
    wire N__39424;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39408;
    wire N__39405;
    wire N__39404;
    wire N__39401;
    wire N__39398;
    wire N__39397;
    wire N__39394;
    wire N__39389;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39315;
    wire N__39314;
    wire N__39309;
    wire N__39308;
    wire N__39307;
    wire N__39304;
    wire N__39299;
    wire N__39294;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39240;
    wire N__39237;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39224;
    wire N__39219;
    wire N__39216;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39204;
    wire N__39203;
    wire N__39200;
    wire N__39197;
    wire N__39194;
    wire N__39189;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39174;
    wire N__39173;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39159;
    wire N__39156;
    wire N__39155;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39138;
    wire N__39137;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39120;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39098;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39078;
    wire N__39075;
    wire N__39070;
    wire N__39067;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38997;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38925;
    wire N__38922;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38843;
    wire N__38840;
    wire N__38837;
    wire N__38834;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38750;
    wire N__38749;
    wire N__38746;
    wire N__38743;
    wire N__38740;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38720;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38708;
    wire N__38705;
    wire N__38702;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38663;
    wire N__38660;
    wire N__38657;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38631;
    wire N__38628;
    wire N__38627;
    wire N__38624;
    wire N__38621;
    wire N__38616;
    wire N__38615;
    wire N__38614;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38546;
    wire N__38543;
    wire N__38540;
    wire N__38535;
    wire N__38532;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38519;
    wire N__38514;
    wire N__38511;
    wire N__38510;
    wire N__38509;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38501;
    wire N__38498;
    wire N__38495;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38472;
    wire N__38469;
    wire N__38468;
    wire N__38465;
    wire N__38464;
    wire N__38461;
    wire N__38460;
    wire N__38459;
    wire N__38458;
    wire N__38453;
    wire N__38452;
    wire N__38451;
    wire N__38448;
    wire N__38443;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38420;
    wire N__38415;
    wire N__38412;
    wire N__38403;
    wire N__38402;
    wire N__38401;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38381;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38356;
    wire N__38351;
    wire N__38348;
    wire N__38345;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38330;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38312;
    wire N__38311;
    wire N__38308;
    wire N__38303;
    wire N__38298;
    wire N__38295;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38265;
    wire N__38262;
    wire N__38261;
    wire N__38260;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38231;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38190;
    wire N__38187;
    wire N__38186;
    wire N__38183;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38167;
    wire N__38160;
    wire N__38157;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38100;
    wire N__38099;
    wire N__38096;
    wire N__38095;
    wire N__38088;
    wire N__38085;
    wire N__38084;
    wire N__38079;
    wire N__38076;
    wire N__38075;
    wire N__38074;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38062;
    wire N__38059;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38043;
    wire N__38042;
    wire N__38041;
    wire N__38038;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37995;
    wire N__37994;
    wire N__37993;
    wire N__37990;
    wire N__37985;
    wire N__37982;
    wire N__37977;
    wire N__37976;
    wire N__37973;
    wire N__37970;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37946;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37908;
    wire N__37905;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37890;
    wire N__37889;
    wire N__37886;
    wire N__37883;
    wire N__37882;
    wire N__37877;
    wire N__37874;
    wire N__37871;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37859;
    wire N__37858;
    wire N__37857;
    wire N__37856;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37811;
    wire N__37810;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37792;
    wire N__37787;
    wire N__37784;
    wire N__37779;
    wire N__37778;
    wire N__37777;
    wire N__37776;
    wire N__37775;
    wire N__37774;
    wire N__37773;
    wire N__37772;
    wire N__37771;
    wire N__37770;
    wire N__37769;
    wire N__37768;
    wire N__37767;
    wire N__37766;
    wire N__37765;
    wire N__37764;
    wire N__37755;
    wire N__37746;
    wire N__37737;
    wire N__37736;
    wire N__37735;
    wire N__37734;
    wire N__37733;
    wire N__37732;
    wire N__37731;
    wire N__37730;
    wire N__37729;
    wire N__37728;
    wire N__37727;
    wire N__37726;
    wire N__37725;
    wire N__37724;
    wire N__37723;
    wire N__37714;
    wire N__37709;
    wire N__37706;
    wire N__37697;
    wire N__37692;
    wire N__37683;
    wire N__37674;
    wire N__37669;
    wire N__37666;
    wire N__37653;
    wire N__37650;
    wire N__37649;
    wire N__37648;
    wire N__37645;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37596;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37581;
    wire N__37578;
    wire N__37577;
    wire N__37572;
    wire N__37571;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37557;
    wire N__37554;
    wire N__37553;
    wire N__37548;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37533;
    wire N__37530;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37518;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37503;
    wire N__37500;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37488;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37473;
    wire N__37470;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37443;
    wire N__37440;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37432;
    wire N__37429;
    wire N__37426;
    wire N__37423;
    wire N__37420;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37392;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37384;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37368;
    wire N__37365;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37357;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37341;
    wire N__37338;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37326;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37311;
    wire N__37308;
    wire N__37307;
    wire N__37306;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37290;
    wire N__37287;
    wire N__37286;
    wire N__37281;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37271;
    wire N__37266;
    wire N__37263;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37251;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37236;
    wire N__37233;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37221;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37206;
    wire N__37203;
    wire N__37202;
    wire N__37199;
    wire N__37196;
    wire N__37195;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37146;
    wire N__37143;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37135;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37119;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37111;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37095;
    wire N__37092;
    wire N__37091;
    wire N__37088;
    wire N__37085;
    wire N__37080;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37065;
    wire N__37062;
    wire N__37061;
    wire N__37056;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37041;
    wire N__37038;
    wire N__37037;
    wire N__37032;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37017;
    wire N__37014;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37002;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36987;
    wire N__36984;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36972;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36957;
    wire N__36954;
    wire N__36953;
    wire N__36950;
    wire N__36947;
    wire N__36944;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36924;
    wire N__36921;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36885;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36794;
    wire N__36791;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36774;
    wire N__36773;
    wire N__36770;
    wire N__36769;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36753;
    wire N__36750;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36701;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36648;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36593;
    wire N__36590;
    wire N__36587;
    wire N__36584;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36441;
    wire N__36440;
    wire N__36435;
    wire N__36434;
    wire N__36433;
    wire N__36432;
    wire N__36431;
    wire N__36430;
    wire N__36427;
    wire N__36416;
    wire N__36415;
    wire N__36410;
    wire N__36407;
    wire N__36402;
    wire N__36399;
    wire N__36398;
    wire N__36397;
    wire N__36392;
    wire N__36389;
    wire N__36388;
    wire N__36387;
    wire N__36384;
    wire N__36377;
    wire N__36372;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36353;
    wire N__36350;
    wire N__36349;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36261;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36195;
    wire N__36192;
    wire N__36191;
    wire N__36188;
    wire N__36185;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36149;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36131;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36116;
    wire N__36115;
    wire N__36112;
    wire N__36111;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36096;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36069;
    wire N__36066;
    wire N__36065;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36048;
    wire N__36045;
    wire N__36044;
    wire N__36041;
    wire N__36040;
    wire N__36037;
    wire N__36036;
    wire N__36033;
    wire N__36026;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35982;
    wire N__35979;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35949;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35927;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35907;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35899;
    wire N__35898;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35862;
    wire N__35859;
    wire N__35858;
    wire N__35853;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35841;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35823;
    wire N__35820;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35799;
    wire N__35796;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35788;
    wire N__35787;
    wire N__35784;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35711;
    wire N__35706;
    wire N__35703;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35684;
    wire N__35681;
    wire N__35678;
    wire N__35673;
    wire N__35672;
    wire N__35671;
    wire N__35668;
    wire N__35663;
    wire N__35660;
    wire N__35655;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35556;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35394;
    wire N__35391;
    wire N__35388;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35378;
    wire N__35375;
    wire N__35374;
    wire N__35371;
    wire N__35370;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35295;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35226;
    wire N__35223;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34971;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34915;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34899;
    wire N__34896;
    wire N__34895;
    wire N__34894;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34878;
    wire N__34875;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34860;
    wire N__34857;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34850;
    wire N__34849;
    wire N__34848;
    wire N__34847;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34838;
    wire N__34837;
    wire N__34836;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34821;
    wire N__34812;
    wire N__34803;
    wire N__34794;
    wire N__34785;
    wire N__34776;
    wire N__34775;
    wire N__34774;
    wire N__34765;
    wire N__34760;
    wire N__34751;
    wire N__34746;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34701;
    wire N__34700;
    wire N__34697;
    wire N__34696;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34675;
    wire N__34672;
    wire N__34667;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34653;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34619;
    wire N__34618;
    wire N__34615;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34593;
    wire N__34590;
    wire N__34589;
    wire N__34588;
    wire N__34587;
    wire N__34586;
    wire N__34585;
    wire N__34584;
    wire N__34583;
    wire N__34582;
    wire N__34581;
    wire N__34580;
    wire N__34579;
    wire N__34578;
    wire N__34577;
    wire N__34576;
    wire N__34575;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34483;
    wire N__34482;
    wire N__34481;
    wire N__34480;
    wire N__34479;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34465;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34449;
    wire N__34442;
    wire N__34433;
    wire N__34424;
    wire N__34415;
    wire N__34412;
    wire N__34405;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34375;
    wire N__34374;
    wire N__34373;
    wire N__34372;
    wire N__34371;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34356;
    wire N__34353;
    wire N__34348;
    wire N__34343;
    wire N__34338;
    wire N__34331;
    wire N__34324;
    wire N__34315;
    wire N__34312;
    wire N__34305;
    wire N__34296;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34290;
    wire N__34287;
    wire N__34280;
    wire N__34269;
    wire N__34262;
    wire N__34259;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34216;
    wire N__34209;
    wire N__34206;
    wire N__34205;
    wire N__34202;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34179;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34145;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34122;
    wire N__34119;
    wire N__34118;
    wire N__34113;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34098;
    wire N__34095;
    wire N__34094;
    wire N__34093;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34077;
    wire N__34074;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34062;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34047;
    wire N__34044;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34036;
    wire N__34031;
    wire N__34028;
    wire N__34025;
    wire N__34020;
    wire N__34017;
    wire N__34016;
    wire N__34015;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__33999;
    wire N__33996;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33974;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33962;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33902;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33865;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33849;
    wire N__33846;
    wire N__33845;
    wire N__33844;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33828;
    wire N__33825;
    wire N__33824;
    wire N__33823;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33807;
    wire N__33804;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33796;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33780;
    wire N__33777;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33765;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33750;
    wire N__33747;
    wire N__33746;
    wire N__33741;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33719;
    wire N__33716;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33699;
    wire N__33696;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33669;
    wire N__33666;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33652;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33636;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33625;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33609;
    wire N__33606;
    wire N__33605;
    wire N__33604;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33588;
    wire N__33585;
    wire N__33584;
    wire N__33583;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33567;
    wire N__33564;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33556;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33533;
    wire N__33530;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33507;
    wire N__33504;
    wire N__33503;
    wire N__33498;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33440;
    wire N__33439;
    wire N__33436;
    wire N__33435;
    wire N__33434;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33405;
    wire N__33402;
    wire N__33397;
    wire N__33394;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33377;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33360;
    wire N__33357;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33303;
    wire N__33302;
    wire N__33299;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33273;
    wire N__33272;
    wire N__33271;
    wire N__33270;
    wire N__33261;
    wire N__33258;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33250;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33236;
    wire N__33231;
    wire N__33228;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33204;
    wire N__33201;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33185;
    wire N__33182;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33128;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33110;
    wire N__33105;
    wire N__33102;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33068;
    wire N__33063;
    wire N__33062;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33047;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33008;
    wire N__33007;
    wire N__33004;
    wire N__32999;
    wire N__32994;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32982;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32967;
    wire N__32966;
    wire N__32965;
    wire N__32964;
    wire N__32963;
    wire N__32962;
    wire N__32961;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32932;
    wire N__32927;
    wire N__32924;
    wire N__32923;
    wire N__32918;
    wire N__32915;
    wire N__32910;
    wire N__32907;
    wire N__32906;
    wire N__32903;
    wire N__32900;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32889;
    wire N__32886;
    wire N__32881;
    wire N__32878;
    wire N__32871;
    wire N__32868;
    wire N__32867;
    wire N__32864;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32831;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32819;
    wire N__32818;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32787;
    wire N__32784;
    wire N__32783;
    wire N__32780;
    wire N__32779;
    wire N__32772;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32760;
    wire N__32757;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32749;
    wire N__32746;
    wire N__32741;
    wire N__32740;
    wire N__32735;
    wire N__32732;
    wire N__32727;
    wire N__32724;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32713;
    wire N__32708;
    wire N__32707;
    wire N__32704;
    wire N__32701;
    wire N__32698;
    wire N__32691;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32657;
    wire N__32652;
    wire N__32649;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32630;
    wire N__32627;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32617;
    wire N__32610;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32591;
    wire N__32588;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32571;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32550;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32522;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32511;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32495;
    wire N__32492;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32480;
    wire N__32477;
    wire N__32474;
    wire N__32473;
    wire N__32470;
    wire N__32465;
    wire N__32464;
    wire N__32459;
    wire N__32456;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32432;
    wire N__32429;
    wire N__32428;
    wire N__32423;
    wire N__32420;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32394;
    wire N__32391;
    wire N__32386;
    wire N__32383;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32369;
    wire N__32366;
    wire N__32363;
    wire N__32358;
    wire N__32357;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32340;
    wire N__32337;
    wire N__32336;
    wire N__32333;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32313;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32295;
    wire N__32292;
    wire N__32291;
    wire N__32288;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32268;
    wire N__32265;
    wire N__32260;
    wire N__32257;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32243;
    wire N__32240;
    wire N__32237;
    wire N__32236;
    wire N__32231;
    wire N__32228;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32187;
    wire N__32180;
    wire N__32177;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32148;
    wire N__32145;
    wire N__32140;
    wire N__32137;
    wire N__32130;
    wire N__32127;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32119;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32105;
    wire N__32102;
    wire N__32101;
    wire N__32096;
    wire N__32093;
    wire N__32088;
    wire N__32085;
    wire N__32084;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32067;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32049;
    wire N__32046;
    wire N__32045;
    wire N__32042;
    wire N__32041;
    wire N__32038;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32022;
    wire N__32019;
    wire N__32014;
    wire N__32011;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31999;
    wire N__31998;
    wire N__31997;
    wire N__31996;
    wire N__31993;
    wire N__31988;
    wire N__31983;
    wire N__31980;
    wire N__31979;
    wire N__31972;
    wire N__31971;
    wire N__31968;
    wire N__31967;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31949;
    wire N__31938;
    wire N__31937;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31896;
    wire N__31895;
    wire N__31892;
    wire N__31891;
    wire N__31890;
    wire N__31887;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31881;
    wire N__31880;
    wire N__31879;
    wire N__31878;
    wire N__31877;
    wire N__31876;
    wire N__31875;
    wire N__31870;
    wire N__31863;
    wire N__31856;
    wire N__31847;
    wire N__31838;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31814;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31793;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31760;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31743;
    wire N__31740;
    wire N__31739;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31726;
    wire N__31723;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31699;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31658;
    wire N__31657;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31634;
    wire N__31633;
    wire N__31630;
    wire N__31625;
    wire N__31624;
    wire N__31619;
    wire N__31616;
    wire N__31611;
    wire N__31608;
    wire N__31607;
    wire N__31604;
    wire N__31601;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31562;
    wire N__31559;
    wire N__31556;
    wire N__31551;
    wire N__31550;
    wire N__31549;
    wire N__31546;
    wire N__31541;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31481;
    wire N__31480;
    wire N__31479;
    wire N__31478;
    wire N__31471;
    wire N__31466;
    wire N__31465;
    wire N__31464;
    wire N__31463;
    wire N__31462;
    wire N__31461;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31442;
    wire N__31439;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31187;
    wire N__31186;
    wire N__31183;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31171;
    wire N__31168;
    wire N__31161;
    wire N__31160;
    wire N__31159;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31147;
    wire N__31144;
    wire N__31137;
    wire N__31136;
    wire N__31135;
    wire N__31132;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31094;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31077;
    wire N__31076;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30948;
    wire N__30947;
    wire N__30946;
    wire N__30945;
    wire N__30944;
    wire N__30943;
    wire N__30942;
    wire N__30939;
    wire N__30932;
    wire N__30927;
    wire N__30926;
    wire N__30925;
    wire N__30924;
    wire N__30923;
    wire N__30922;
    wire N__30921;
    wire N__30920;
    wire N__30919;
    wire N__30918;
    wire N__30917;
    wire N__30916;
    wire N__30915;
    wire N__30912;
    wire N__30911;
    wire N__30910;
    wire N__30909;
    wire N__30908;
    wire N__30907;
    wire N__30904;
    wire N__30899;
    wire N__30884;
    wire N__30871;
    wire N__30860;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30846;
    wire N__30843;
    wire N__30834;
    wire N__30831;
    wire N__30830;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30812;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30692;
    wire N__30691;
    wire N__30690;
    wire N__30689;
    wire N__30688;
    wire N__30687;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30679;
    wire N__30678;
    wire N__30677;
    wire N__30676;
    wire N__30675;
    wire N__30674;
    wire N__30673;
    wire N__30672;
    wire N__30671;
    wire N__30670;
    wire N__30669;
    wire N__30668;
    wire N__30667;
    wire N__30666;
    wire N__30665;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30625;
    wire N__30624;
    wire N__30623;
    wire N__30622;
    wire N__30621;
    wire N__30620;
    wire N__30619;
    wire N__30616;
    wire N__30615;
    wire N__30614;
    wire N__30611;
    wire N__30610;
    wire N__30607;
    wire N__30606;
    wire N__30605;
    wire N__30604;
    wire N__30603;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30597;
    wire N__30596;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30567;
    wire N__30566;
    wire N__30563;
    wire N__30560;
    wire N__30555;
    wire N__30548;
    wire N__30545;
    wire N__30538;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30493;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30475;
    wire N__30472;
    wire N__30471;
    wire N__30470;
    wire N__30469;
    wire N__30468;
    wire N__30467;
    wire N__30466;
    wire N__30465;
    wire N__30464;
    wire N__30461;
    wire N__30460;
    wire N__30459;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30448;
    wire N__30445;
    wire N__30444;
    wire N__30443;
    wire N__30442;
    wire N__30441;
    wire N__30440;
    wire N__30439;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30435;
    wire N__30434;
    wire N__30433;
    wire N__30432;
    wire N__30431;
    wire N__30430;
    wire N__30429;
    wire N__30428;
    wire N__30427;
    wire N__30426;
    wire N__30425;
    wire N__30424;
    wire N__30421;
    wire N__30412;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30393;
    wire N__30390;
    wire N__30375;
    wire N__30366;
    wire N__30359;
    wire N__30354;
    wire N__30351;
    wire N__30350;
    wire N__30349;
    wire N__30348;
    wire N__30347;
    wire N__30346;
    wire N__30343;
    wire N__30338;
    wire N__30335;
    wire N__30334;
    wire N__30333;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30316;
    wire N__30309;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30286;
    wire N__30285;
    wire N__30284;
    wire N__30283;
    wire N__30282;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30278;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30274;
    wire N__30273;
    wire N__30272;
    wire N__30269;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30186;
    wire N__30183;
    wire N__30176;
    wire N__30171;
    wire N__30164;
    wire N__30157;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30145;
    wire N__30142;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30104;
    wire N__30099;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30036;
    wire N__30033;
    wire N__30024;
    wire N__30015;
    wire N__30006;
    wire N__29997;
    wire N__29988;
    wire N__29981;
    wire N__29974;
    wire N__29969;
    wire N__29960;
    wire N__29953;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29937;
    wire N__29930;
    wire N__29921;
    wire N__29912;
    wire N__29903;
    wire N__29898;
    wire N__29879;
    wire N__29870;
    wire N__29847;
    wire N__29846;
    wire N__29845;
    wire N__29844;
    wire N__29843;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29837;
    wire N__29836;
    wire N__29835;
    wire N__29834;
    wire N__29833;
    wire N__29832;
    wire N__29829;
    wire N__29828;
    wire N__29825;
    wire N__29824;
    wire N__29823;
    wire N__29822;
    wire N__29821;
    wire N__29820;
    wire N__29819;
    wire N__29818;
    wire N__29817;
    wire N__29816;
    wire N__29815;
    wire N__29814;
    wire N__29813;
    wire N__29812;
    wire N__29811;
    wire N__29810;
    wire N__29809;
    wire N__29808;
    wire N__29807;
    wire N__29804;
    wire N__29803;
    wire N__29802;
    wire N__29801;
    wire N__29800;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29784;
    wire N__29783;
    wire N__29782;
    wire N__29777;
    wire N__29768;
    wire N__29767;
    wire N__29764;
    wire N__29761;
    wire N__29756;
    wire N__29747;
    wire N__29740;
    wire N__29737;
    wire N__29736;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29722;
    wire N__29719;
    wire N__29710;
    wire N__29709;
    wire N__29708;
    wire N__29707;
    wire N__29706;
    wire N__29705;
    wire N__29704;
    wire N__29703;
    wire N__29702;
    wire N__29701;
    wire N__29700;
    wire N__29699;
    wire N__29698;
    wire N__29697;
    wire N__29696;
    wire N__29693;
    wire N__29692;
    wire N__29691;
    wire N__29690;
    wire N__29687;
    wire N__29682;
    wire N__29675;
    wire N__29670;
    wire N__29665;
    wire N__29662;
    wire N__29651;
    wire N__29648;
    wire N__29639;
    wire N__29634;
    wire N__29631;
    wire N__29630;
    wire N__29625;
    wire N__29618;
    wire N__29609;
    wire N__29600;
    wire N__29595;
    wire N__29592;
    wire N__29591;
    wire N__29588;
    wire N__29585;
    wire N__29582;
    wire N__29581;
    wire N__29580;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29563;
    wire N__29550;
    wire N__29547;
    wire N__29536;
    wire N__29535;
    wire N__29534;
    wire N__29529;
    wire N__29524;
    wire N__29521;
    wire N__29516;
    wire N__29513;
    wire N__29504;
    wire N__29501;
    wire N__29496;
    wire N__29491;
    wire N__29484;
    wire N__29481;
    wire N__29466;
    wire N__29465;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29455;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29392;
    wire N__29387;
    wire N__29384;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29373;
    wire N__29370;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29330;
    wire N__29327;
    wire N__29322;
    wire N__29321;
    wire N__29320;
    wire N__29317;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29281;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29252;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29212;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29200;
    wire N__29193;
    wire N__29190;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29182;
    wire N__29181;
    wire N__29176;
    wire N__29171;
    wire N__29168;
    wire N__29165;
    wire N__29160;
    wire N__29159;
    wire N__29158;
    wire N__29153;
    wire N__29152;
    wire N__29149;
    wire N__29148;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29122;
    wire N__29115;
    wire N__29112;
    wire N__29111;
    wire N__29110;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29100;
    wire N__29099;
    wire N__29098;
    wire N__29095;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29087;
    wire N__29086;
    wire N__29085;
    wire N__29084;
    wire N__29083;
    wire N__29068;
    wire N__29065;
    wire N__29060;
    wire N__29059;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29039;
    wire N__29038;
    wire N__29037;
    wire N__29034;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29010;
    wire N__29003;
    wire N__28998;
    wire N__28993;
    wire N__28980;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28968;
    wire N__28967;
    wire N__28966;
    wire N__28965;
    wire N__28964;
    wire N__28963;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28946;
    wire N__28945;
    wire N__28944;
    wire N__28943;
    wire N__28942;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28936;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28928;
    wire N__28927;
    wire N__28924;
    wire N__28913;
    wire N__28906;
    wire N__28891;
    wire N__28888;
    wire N__28887;
    wire N__28884;
    wire N__28883;
    wire N__28878;
    wire N__28875;
    wire N__28870;
    wire N__28867;
    wire N__28866;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28850;
    wire N__28847;
    wire N__28836;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28828;
    wire N__28827;
    wire N__28826;
    wire N__28825;
    wire N__28824;
    wire N__28823;
    wire N__28822;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28815;
    wire N__28814;
    wire N__28797;
    wire N__28790;
    wire N__28785;
    wire N__28770;
    wire N__28769;
    wire N__28768;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28751;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28732;
    wire N__28729;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28703;
    wire N__28700;
    wire N__28699;
    wire N__28698;
    wire N__28695;
    wire N__28694;
    wire N__28693;
    wire N__28692;
    wire N__28691;
    wire N__28688;
    wire N__28687;
    wire N__28686;
    wire N__28677;
    wire N__28672;
    wire N__28671;
    wire N__28668;
    wire N__28667;
    wire N__28664;
    wire N__28659;
    wire N__28654;
    wire N__28647;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28619;
    wire N__28616;
    wire N__28613;
    wire N__28608;
    wire N__28605;
    wire N__28604;
    wire N__28599;
    wire N__28598;
    wire N__28597;
    wire N__28594;
    wire N__28589;
    wire N__28584;
    wire N__28583;
    wire N__28578;
    wire N__28577;
    wire N__28574;
    wire N__28571;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28506;
    wire N__28505;
    wire N__28502;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28485;
    wire N__28482;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28474;
    wire N__28469;
    wire N__28466;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28426;
    wire N__28421;
    wire N__28418;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28400;
    wire N__28399;
    wire N__28396;
    wire N__28391;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28363;
    wire N__28358;
    wire N__28355;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28330;
    wire N__28325;
    wire N__28322;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28205;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28142;
    wire N__28141;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28111;
    wire N__28106;
    wire N__28103;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28075;
    wire N__28070;
    wire N__28067;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28039;
    wire N__28034;
    wire N__28031;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27998;
    wire N__27997;
    wire N__27992;
    wire N__27989;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27974;
    wire N__27973;
    wire N__27970;
    wire N__27965;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27943;
    wire N__27938;
    wire N__27935;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27882;
    wire N__27881;
    wire N__27878;
    wire N__27875;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27863;
    wire N__27862;
    wire N__27859;
    wire N__27854;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27836;
    wire N__27831;
    wire N__27828;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27764;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27731;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27696;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27653;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27626;
    wire N__27625;
    wire N__27622;
    wire N__27617;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27602;
    wire N__27601;
    wire N__27598;
    wire N__27593;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27473;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27089;
    wire N__27088;
    wire N__27087;
    wire N__27086;
    wire N__27085;
    wire N__27084;
    wire N__27083;
    wire N__27082;
    wire N__27081;
    wire N__27080;
    wire N__27079;
    wire N__27078;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27054;
    wire N__27041;
    wire N__27038;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27026;
    wire N__27025;
    wire N__27024;
    wire N__27023;
    wire N__27022;
    wire N__27021;
    wire N__27020;
    wire N__27019;
    wire N__27018;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27006;
    wire N__26997;
    wire N__26986;
    wire N__26983;
    wire N__26970;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26696;
    wire N__26695;
    wire N__26694;
    wire N__26691;
    wire N__26684;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26484;
    wire N__26481;
    wire N__26478;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26340;
    wire N__26337;
    wire N__26334;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26315;
    wire N__26312;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26295;
    wire N__26292;
    wire N__26289;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26277;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26256;
    wire N__26253;
    wire N__26250;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25995;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25016;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24945;
    wire N__24942;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24917;
    wire N__24916;
    wire N__24915;
    wire N__24914;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24906;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24884;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24872;
    wire N__24871;
    wire N__24868;
    wire N__24867;
    wire N__24866;
    wire N__24863;
    wire N__24862;
    wire N__24861;
    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24826;
    wire N__24825;
    wire N__24824;
    wire N__24823;
    wire N__24822;
    wire N__24821;
    wire N__24816;
    wire N__24813;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24805;
    wire N__24800;
    wire N__24797;
    wire N__24790;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24775;
    wire N__24774;
    wire N__24771;
    wire N__24770;
    wire N__24767;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24752;
    wire N__24749;
    wire N__24748;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24703;
    wire N__24700;
    wire N__24695;
    wire N__24690;
    wire N__24687;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24664;
    wire N__24661;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24629;
    wire N__24622;
    wire N__24617;
    wire N__24614;
    wire N__24609;
    wire N__24606;
    wire N__24601;
    wire N__24596;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24506;
    wire N__24501;
    wire N__24498;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24456;
    wire N__24453;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24431;
    wire N__24428;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24411;
    wire N__24408;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24267;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24201;
    wire N__24198;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24128;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24096;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24054;
    wire N__24051;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23978;
    wire N__23975;
    wire N__23974;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23953;
    wire N__23950;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23920;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23916;
    wire N__23915;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23907;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23901;
    wire N__23900;
    wire N__23899;
    wire N__23898;
    wire N__23897;
    wire N__23892;
    wire N__23889;
    wire N__23882;
    wire N__23871;
    wire N__23870;
    wire N__23869;
    wire N__23868;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23864;
    wire N__23863;
    wire N__23862;
    wire N__23855;
    wire N__23852;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23834;
    wire N__23827;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23796;
    wire N__23795;
    wire N__23794;
    wire N__23785;
    wire N__23782;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23760;
    wire N__23759;
    wire N__23758;
    wire N__23757;
    wire N__23756;
    wire N__23755;
    wire N__23748;
    wire N__23747;
    wire N__23746;
    wire N__23745;
    wire N__23742;
    wire N__23737;
    wire N__23736;
    wire N__23735;
    wire N__23734;
    wire N__23733;
    wire N__23732;
    wire N__23731;
    wire N__23730;
    wire N__23729;
    wire N__23728;
    wire N__23725;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23702;
    wire N__23691;
    wire N__23690;
    wire N__23689;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23684;
    wire N__23683;
    wire N__23682;
    wire N__23681;
    wire N__23680;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23670;
    wire N__23661;
    wire N__23648;
    wire N__23633;
    wire N__23622;
    wire N__23621;
    wire N__23620;
    wire N__23619;
    wire N__23618;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23611;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23603;
    wire N__23602;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23589;
    wire N__23588;
    wire N__23585;
    wire N__23584;
    wire N__23583;
    wire N__23582;
    wire N__23581;
    wire N__23580;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23566;
    wire N__23565;
    wire N__23558;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23539;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23472;
    wire N__23469;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23449;
    wire N__23440;
    wire N__23437;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23417;
    wire N__23414;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23381;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23361;
    wire N__23358;
    wire N__23357;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23337;
    wire N__23336;
    wire N__23333;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23316;
    wire N__23315;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23274;
    wire N__23273;
    wire N__23270;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23253;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23245;
    wire N__23240;
    wire N__23237;
    wire N__23232;
    wire N__23229;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23221;
    wire N__23216;
    wire N__23213;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23201;
    wire N__23198;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23174;
    wire N__23173;
    wire N__23170;
    wire N__23167;
    wire N__23164;
    wire N__23157;
    wire N__23156;
    wire N__23155;
    wire N__23154;
    wire N__23153;
    wire N__23152;
    wire N__23151;
    wire N__23150;
    wire N__23149;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23133;
    wire N__23124;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23096;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23068;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23051;
    wire N__23050;
    wire N__23045;
    wire N__23042;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22996;
    wire N__22993;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22975;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22958;
    wire N__22957;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22918;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22886;
    wire N__22885;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22852;
    wire N__22851;
    wire N__22848;
    wire N__22843;
    wire N__22840;
    wire N__22833;
    wire N__22830;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22822;
    wire N__22821;
    wire N__22818;
    wire N__22813;
    wire N__22810;
    wire N__22805;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22787;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22773;
    wire N__22770;
    wire N__22765;
    wire N__22762;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22736;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22718;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22681;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22658;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22591;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22571;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22534;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22520;
    wire N__22517;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22492;
    wire N__22485;
    wire N__22482;
    wire N__22481;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22449;
    wire N__22446;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22438;
    wire N__22437;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22416;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22408;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22374;
    wire N__22371;
    wire N__22370;
    wire N__22367;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22278;
    wire N__22275;
    wire N__22270;
    wire N__22267;
    wire N__22262;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22231;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22208;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22196;
    wire N__22193;
    wire N__22192;
    wire N__22189;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22168;
    wire N__22165;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22138;
    wire N__22135;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22111;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22064;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22056;
    wire N__22053;
    wire N__22048;
    wire N__22045;
    wire N__22038;
    wire N__22037;
    wire N__22034;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22017;
    wire N__22016;
    wire N__22015;
    wire N__22014;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21973;
    wire N__21970;
    wire N__21965;
    wire N__21954;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21897;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21885;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21870;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21858;
    wire N__21855;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21843;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21831;
    wire N__21828;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21813;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21783;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21771;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21680;
    wire N__21675;
    wire N__21674;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21617;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21590;
    wire N__21589;
    wire N__21586;
    wire N__21585;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21569;
    wire N__21566;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21542;
    wire N__21541;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21529;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21493;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21467;
    wire N__21464;
    wire N__21463;
    wire N__21462;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21377;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21118;
    wire N__21117;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20873;
    wire N__20870;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20837;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20801;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20768;
    wire N__20765;
    wire N__20762;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20747;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20573;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20540;
    wire N__20537;
    wire N__20536;
    wire N__20535;
    wire N__20534;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20522;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20503;
    wire N__20500;
    wire N__20487;
    wire N__20480;
    wire N__20475;
    wire N__20472;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20423;
    wire N__20422;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20414;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20403;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20347;
    wire N__20340;
    wire N__20339;
    wire N__20338;
    wire N__20337;
    wire N__20336;
    wire N__20335;
    wire N__20334;
    wire N__20331;
    wire N__20330;
    wire N__20329;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20307;
    wire N__20306;
    wire N__20301;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20285;
    wire N__20280;
    wire N__20279;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20275;
    wire N__20274;
    wire N__20271;
    wire N__20270;
    wire N__20269;
    wire N__20264;
    wire N__20263;
    wire N__20262;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20251;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20239;
    wire N__20238;
    wire N__20237;
    wire N__20236;
    wire N__20235;
    wire N__20234;
    wire N__20233;
    wire N__20232;
    wire N__20229;
    wire N__20222;
    wire N__20215;
    wire N__20210;
    wire N__20207;
    wire N__20202;
    wire N__20201;
    wire N__20200;
    wire N__20199;
    wire N__20198;
    wire N__20197;
    wire N__20196;
    wire N__20195;
    wire N__20194;
    wire N__20193;
    wire N__20192;
    wire N__20191;
    wire N__20176;
    wire N__20171;
    wire N__20162;
    wire N__20157;
    wire N__20154;
    wire N__20137;
    wire N__20132;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19959;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19881;
    wire N__19878;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19830;
    wire N__19827;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19815;
    wire N__19812;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19764;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19749;
    wire N__19748;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19725;
    wire N__19722;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19704;
    wire N__19701;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19683;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19665;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19610;
    wire N__19607;
    wire N__19606;
    wire N__19605;
    wire N__19604;
    wire N__19601;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19587;
    wire N__19586;
    wire N__19583;
    wire N__19582;
    wire N__19581;
    wire N__19580;
    wire N__19573;
    wire N__19570;
    wire N__19561;
    wire N__19558;
    wire N__19553;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19530;
    wire N__19527;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19502;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19491;
    wire N__19488;
    wire N__19481;
    wire N__19480;
    wire N__19479;
    wire N__19478;
    wire N__19477;
    wire N__19472;
    wire N__19469;
    wire N__19462;
    wire N__19459;
    wire N__19454;
    wire N__19449;
    wire N__19446;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19364;
    wire N__19359;
    wire N__19356;
    wire N__19355;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19331;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19223;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19205;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19193;
    wire N__19192;
    wire N__19191;
    wire N__19188;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19172;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19157;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19133;
    wire N__19128;
    wire N__19125;
    wire N__19124;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19106;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19094;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19076;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19035;
    wire N__19034;
    wire N__19029;
    wire N__19026;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18884;
    wire N__18883;
    wire N__18882;
    wire N__18881;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18867;
    wire N__18864;
    wire N__18855;
    wire N__18852;
    wire N__18851;
    wire N__18848;
    wire N__18847;
    wire N__18844;
    wire N__18839;
    wire N__18836;
    wire N__18831;
    wire N__18828;
    wire N__18827;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18731;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18681;
    wire N__18680;
    wire N__18677;
    wire N__18676;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18214;
    wire N__18213;
    wire N__18212;
    wire N__18207;
    wire N__18204;
    wire N__18203;
    wire N__18200;
    wire N__18199;
    wire N__18196;
    wire N__18195;
    wire N__18192;
    wire N__18179;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17955;
    wire N__17952;
    wire N__17951;
    wire N__17950;
    wire N__17947;
    wire N__17942;
    wire N__17939;
    wire N__17934;
    wire N__17933;
    wire N__17932;
    wire N__17929;
    wire N__17924;
    wire N__17921;
    wire N__17916;
    wire N__17915;
    wire N__17914;
    wire N__17911;
    wire N__17906;
    wire N__17903;
    wire N__17898;
    wire N__17895;
    wire N__17894;
    wire N__17893;
    wire N__17890;
    wire N__17885;
    wire N__17882;
    wire N__17877;
    wire N__17876;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17856;
    wire N__17853;
    wire N__17852;
    wire N__17851;
    wire N__17848;
    wire N__17843;
    wire N__17840;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ;
    wire pwm_duty_input_6;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire pwm_duty_input_4;
    wire pwm_duty_input_8;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire bfn_1_12_0_;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_1_13_0_;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire bfn_1_16_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire un7_start_stop_0_a3;
    wire N_34_i_i;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire bfn_2_7_0_;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire bfn_2_8_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_94_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_120 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.N_118_cascade_ ;
    wire pwm_duty_input_9;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_2_13_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_2_14_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire bfn_2_15_0_;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire bfn_2_16_0_;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.N_16 ;
    wire N_19_1;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_3_10_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_3_11_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire bfn_3_18_0_;
    wire un5_counter_cry_1;
    wire un5_counter_cry_2;
    wire un5_counter_cry_3;
    wire un5_counter_cry_4;
    wire un5_counter_cry_5;
    wire un5_counter_cry_6;
    wire un5_counter_cry_7;
    wire un5_counter_cry_8;
    wire bfn_3_19_0_;
    wire un5_counter_cry_9;
    wire un5_counter_cry_10;
    wire un5_counter_cry_11;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_4_6_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_4_7_0_;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \current_shift_inst.PI_CTRL.N_170_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.N_168 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire bfn_4_13_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire bfn_4_14_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire bfn_4_15_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire bfn_4_16_0_;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire counterZ0Z_11;
    wire counterZ0Z_6;
    wire counterZ0Z_12;
    wire counterZ0Z_10;
    wire \current_shift_inst.PI_CTRL.un2_counterZ0Z_1_cascade_ ;
    wire counterZ0Z_8;
    wire counterZ0Z_7;
    wire counterZ0Z_9;
    wire counterZ0Z_5;
    wire \current_shift_inst.PI_CTRL.un2_counterZ0Z_8 ;
    wire counterZ0Z_2;
    wire counterZ0Z_3;
    wire counterZ0Z_4;
    wire \current_shift_inst.PI_CTRL.un2_counterZ0Z_7 ;
    wire counterZ0Z_1;
    wire counterZ0Z_0;
    wire \current_shift_inst.PI_CTRL.un2_counterZ0 ;
    wire clk_10khz_i;
    wire bfn_5_6_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_5_7_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.N_167 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.N_171_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_170 ;
    wire \current_shift_inst.PI_CTRL.N_171 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire il_max_comp2_c;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.control_inputZ0Z_0 ;
    wire bfn_7_13_0_;
    wire \current_shift_inst.control_inputZ0Z_1 ;
    wire \current_shift_inst.control_input_1_cry_0 ;
    wire \current_shift_inst.control_inputZ0Z_2 ;
    wire \current_shift_inst.control_input_1_cry_1 ;
    wire \current_shift_inst.control_inputZ0Z_3 ;
    wire \current_shift_inst.control_input_1_cry_2 ;
    wire \current_shift_inst.control_inputZ0Z_4 ;
    wire \current_shift_inst.control_input_1_cry_3 ;
    wire \current_shift_inst.control_inputZ0Z_5 ;
    wire \current_shift_inst.control_input_1_cry_4 ;
    wire \current_shift_inst.control_inputZ0Z_6 ;
    wire \current_shift_inst.control_input_1_cry_5 ;
    wire \current_shift_inst.control_inputZ0Z_7 ;
    wire \current_shift_inst.control_input_1_cry_6 ;
    wire \current_shift_inst.control_input_1_cry_7 ;
    wire \current_shift_inst.control_inputZ0Z_8 ;
    wire bfn_7_14_0_;
    wire \current_shift_inst.control_inputZ0Z_9 ;
    wire \current_shift_inst.control_input_1_cry_8 ;
    wire \current_shift_inst.control_inputZ0Z_10 ;
    wire \current_shift_inst.control_input_1_cry_9 ;
    wire \current_shift_inst.control_inputZ0Z_11 ;
    wire \current_shift_inst.control_input_1_cry_10 ;
    wire \current_shift_inst.control_inputZ0Z_12 ;
    wire \current_shift_inst.control_input_1_cry_11 ;
    wire \current_shift_inst.control_inputZ0Z_13 ;
    wire \current_shift_inst.control_input_1_cry_12 ;
    wire \current_shift_inst.control_inputZ0Z_14 ;
    wire \current_shift_inst.control_input_1_cry_13 ;
    wire \current_shift_inst.control_inputZ0Z_15 ;
    wire \current_shift_inst.control_input_1_cry_14 ;
    wire \current_shift_inst.control_input_1_cry_15 ;
    wire \current_shift_inst.control_inputZ0Z_16 ;
    wire bfn_7_15_0_;
    wire \current_shift_inst.control_inputZ0Z_17 ;
    wire \current_shift_inst.control_input_1_cry_16 ;
    wire \current_shift_inst.control_inputZ0Z_18 ;
    wire \current_shift_inst.control_input_1_cry_17 ;
    wire \current_shift_inst.control_inputZ0Z_19 ;
    wire \current_shift_inst.control_input_1_cry_18 ;
    wire \current_shift_inst.control_inputZ0Z_20 ;
    wire \current_shift_inst.control_input_1_cry_19 ;
    wire \current_shift_inst.control_inputZ0Z_21 ;
    wire \current_shift_inst.control_input_1_cry_20 ;
    wire \current_shift_inst.control_inputZ0Z_22 ;
    wire \current_shift_inst.control_input_1_cry_21 ;
    wire \current_shift_inst.control_inputZ0Z_23 ;
    wire \current_shift_inst.control_input_1_cry_22 ;
    wire \current_shift_inst.control_input_1_cry_23 ;
    wire \current_shift_inst.control_inputZ0Z_24 ;
    wire bfn_7_16_0_;
    wire \current_shift_inst.control_input_1_cry_24 ;
    wire \current_shift_inst.control_inputZ0Z_25 ;
    wire N_748_g;
    wire \current_shift_inst.control_input_1_axb_23 ;
    wire il_max_comp1_c;
    wire il_min_comp2_c;
    wire il_min_comp2_D1;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire bfn_8_11_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_8_12_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire bfn_8_13_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ;
    wire \current_shift_inst.control_input_1_axb_22 ;
    wire \current_shift_inst.control_input_1_axb_21 ;
    wire \current_shift_inst.control_input_1_axb_3 ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire \current_shift_inst.control_input_1_axb_2 ;
    wire \current_shift_inst.control_input_1_axb_6 ;
    wire \current_shift_inst.control_input_1_axb_5 ;
    wire \current_shift_inst.control_input_1_axb_14 ;
    wire \current_shift_inst.control_input_1_axb_13 ;
    wire \current_shift_inst.control_input_1_axb_12 ;
    wire \current_shift_inst.control_input_1_axb_15 ;
    wire \current_shift_inst.control_input_1_axb_10 ;
    wire \current_shift_inst.control_input_1_axb_16 ;
    wire \current_shift_inst.control_input_1_axb_11 ;
    wire \current_shift_inst.control_input_1_axb_8 ;
    wire \current_shift_inst.control_input_1_axb_20 ;
    wire \current_shift_inst.control_input_1_axb_0 ;
    wire \current_shift_inst.control_input_1_axb_18 ;
    wire \current_shift_inst.control_input_1_axb_19 ;
    wire \current_shift_inst.control_input_1_axb_24 ;
    wire \current_shift_inst.control_input_1_axb_9 ;
    wire \current_shift_inst.control_input_1_axb_1 ;
    wire \current_shift_inst.control_input_1_axb_17 ;
    wire \current_shift_inst.control_input_1_axb_4 ;
    wire \current_shift_inst.control_input_1_axb_7 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_1_axb_25 ;
    wire s4_phy_c;
    wire il_max_comp1_D1;
    wire il_max_comp2_D1;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ;
    wire bfn_9_15_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_9_16_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_9_22_0_;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire s3_phy_c;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_10_11_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_10_12_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_17 ;
    wire bfn_10_13_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.N_1819_i ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire il_max_comp2_D2;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_11_14_0_;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_0_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_463_i ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_257 ;
    wire \phase_controller_inst1.stoper_tr.N_257_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_240 ;
    wire start_stop_c;
    wire \phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \phase_controller_inst2.stoper_tr.time_passed11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire state_ns_i_a3_1;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_185_i ;
    wire \delay_measurement_inst.prev_tr_sigZ0 ;
    wire \delay_measurement_inst.tr_stateZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hc_RNO_0_0 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_13_8_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_13_9_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_17 ;
    wire bfn_13_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire measured_delay_tr_15;
    wire measured_delay_tr_14;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ;
    wire \delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14 ;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_13_15_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_13_16_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_13_17_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_13_18_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_185_i_g ;
    wire s1_phy_c;
    wire delay_tr_input_c;
    wire delay_tr_d1;
    wire delay_tr_d2;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ;
    wire pwm_duty_input_1;
    wire pwm_duty_input_0;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \phase_controller_inst1.stoper_tr.time_passed11_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ;
    wire \delay_measurement_inst.N_360_cascade_ ;
    wire measured_delay_tr_9;
    wire \delay_measurement_inst.N_354_cascade_ ;
    wire measured_delay_tr_10;
    wire measured_delay_tr_11;
    wire measured_delay_tr_12;
    wire \delay_measurement_inst.N_354 ;
    wire measured_delay_tr_13;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_14_13_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_186_i ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_14_19_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire bfn_14_20_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_16 ;
    wire bfn_14_21_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ;
    wire bfn_14_25_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_14_26_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_14_27_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_14_28_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire il_min_comp1_D1;
    wire \phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_15_8_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ;
    wire bfn_15_9_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ;
    wire bfn_15_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31_cascade_ ;
    wire measured_delay_tr_6;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0 ;
    wire \delay_measurement_inst.N_381_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_376 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_ ;
    wire \delay_measurement_inst.N_498_cascade_ ;
    wire \delay_measurement_inst.N_381 ;
    wire \delay_measurement_inst.N_384 ;
    wire \delay_measurement_inst.N_384_cascade_ ;
    wire measured_delay_tr_4;
    wire measured_delay_tr_5;
    wire measured_delay_tr_7;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31 ;
    wire measured_delay_tr_8;
    wire measured_delay_tr_3;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_hc_RNOZ0Z_0_cascade_ ;
    wire il_max_comp1_D2;
    wire state_3;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire s2_phy_c;
    wire measured_delay_tr_1;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i ;
    wire \delay_measurement_inst.delay_tr_reg_5_tz_1 ;
    wire measured_delay_tr_2;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_15_17_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire bfn_15_18_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire bfn_15_19_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_15_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_15_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_15_24_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_15_25_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_461_i_g ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_462_i ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0 ;
    wire \phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_ ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.stoper_tr.time_passed11 ;
    wire \phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire measured_delay_tr_16;
    wire measured_delay_tr_19;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ;
    wire \delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_6 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \delay_measurement_inst.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ;
    wire \delay_measurement_inst.delay_tr_timer.N_373_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ;
    wire \delay_measurement_inst.elapsed_time_tr_3 ;
    wire bfn_16_11_0_;
    wire \delay_measurement_inst.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_reg3lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_reg3lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.elapsed_time_tr_11 ;
    wire bfn_16_12_0_;
    wire \delay_measurement_inst.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_reg3lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_reg3lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.elapsed_time_tr_19 ;
    wire bfn_16_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_16_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0Z0Z_3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_316_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un2_startlt31_5_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.N_406 ;
    wire \phase_controller_inst1.stoper_hc.N_406_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.time_passed11 ;
    wire \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_7_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2Z0Z_18 ;
    wire \delay_measurement_inst.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.elapsed_time_hc_10 ;
    wire measured_delay_hc_24;
    wire measured_delay_hc_23;
    wire measured_delay_hc_22;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7Z0Z_19_cascade_ ;
    wire \delay_measurement_inst.delay_hc_reg3lto14 ;
    wire \delay_measurement_inst.delay_hc_reg3lto9 ;
    wire \delay_measurement_inst.delay_hc_timer.N_299_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_2_6 ;
    wire \delay_measurement_inst.N_332_cascade_ ;
    wire \delay_measurement_inst.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.N_318_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_440 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_0_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_328_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_4 ;
    wire \delay_measurement_inst.delay_hc_timer.N_318_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_331 ;
    wire \delay_measurement_inst.delay_hc_timer.N_328 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_319 ;
    wire \delay_measurement_inst.N_318_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_6_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_7_6 ;
    wire measured_delay_hc_21;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0Z0Z_19 ;
    wire \delay_measurement_inst.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.N_408 ;
    wire measured_delay_hc_26;
    wire \delay_measurement_inst.elapsed_time_hc_17 ;
    wire measured_delay_hc_20;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_461_i ;
    wire delay_hc_input_c;
    wire delay_hc_d1;
    wire bfn_17_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_17_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_464_i ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ;
    wire \phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ;
    wire \delay_measurement_inst.hc_stateZ0Z_0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa_cascade_ ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire delay_hc_d2;
    wire \delay_measurement_inst.prev_hc_sigZ0 ;
    wire measured_delay_hc_8;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1 ;
    wire measured_delay_hc_7;
    wire measured_delay_hc_5;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3Z0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.N_388 ;
    wire \phase_controller_inst1.stoper_hc.N_405_cascade_ ;
    wire measured_delay_hc_4;
    wire measured_delay_hc_10;
    wire measured_delay_hc_11;
    wire measured_delay_hc_12;
    wire measured_delay_hc_13;
    wire \phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.N_459 ;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3 ;
    wire measured_delay_hc_3;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3_cascade_ ;
    wire measured_delay_hc_14;
    wire \phase_controller_inst1.stoper_hc.N_405 ;
    wire measured_delay_hc_9;
    wire measured_delay_hc_30;
    wire \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6Z0Z_19 ;
    wire measured_delay_hc_6;
    wire measured_delay_hc_29;
    wire measured_delay_hc_27;
    wire measured_delay_hc_28;
    wire measured_delay_hc_0;
    wire \delay_measurement_inst.elapsed_time_hc_19 ;
    wire measured_delay_hc_19;
    wire \delay_measurement_inst.elapsed_time_hc_16 ;
    wire measured_delay_hc_1;
    wire \delay_measurement_inst.elapsed_time_hc_18 ;
    wire measured_delay_hc_18;
    wire \delay_measurement_inst.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.elapsed_time_hc_3 ;
    wire \delay_measurement_inst.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_3 ;
    wire \delay_measurement_inst.delay_hc_reg3lto6 ;
    wire \delay_measurement_inst.N_332 ;
    wire \delay_measurement_inst.N_318 ;
    wire \delay_measurement_inst.N_295 ;
    wire \delay_measurement_inst.delay_hc_reg3lto15 ;
    wire measured_delay_hc_15;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_463_i_g ;
    wire \delay_measurement_inst.elapsed_time_tr_17 ;
    wire measured_delay_tr_17;
    wire \delay_measurement_inst.N_498 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.elapsed_time_tr_18 ;
    wire measured_delay_tr_18;
    wire \delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ;
    wire red_c_i;
    wire \phase_controller_inst2.stoper_hc.time_passed11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ;
    wire bfn_18_13_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ;
    wire bfn_18_14_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ;
    wire bfn_18_15_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ;
    wire \phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ;
    wire bfn_18_17_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire bfn_18_18_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_16 ;
    wire bfn_18_19_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.N_453 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire measured_delay_hc_16;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.N_449 ;
    wire measured_delay_hc_31;
    wire measured_delay_hc_17;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ;
    wire measured_delay_hc_25;
    wire \delay_measurement_inst.N_312 ;
    wire \delay_measurement_inst.elapsed_time_hc_2 ;
    wire \delay_measurement_inst.N_298 ;
    wire measured_delay_hc_2;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__18576),
            .RESETB(N__42506),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__34374),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__34367),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__20197,N__20238,N__20195,N__20237,N__20196,N__20236,N__20198,N__20233,N__20191,N__20232,N__20192,N__20234,N__20193,N__20235,N__20194}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__34373,N__34370,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__34368,N__34372,N__34369,N__34371}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__34565),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__34558),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__20261,N__20278,N__20262,N__20279,N__20263,N__18851,N__17877,N__17934,N__17952,N__17916,N__17898,N__17853,N__33170,N__33227,N__33200}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__34564,N__34561,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__34559,N__34563,N__34560,N__34562}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__47200),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__47202),
            .DIN(N__47201),
            .DOUT(N__47200),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__47202),
            .PADOUT(N__47201),
            .PADIN(N__47200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__47191),
            .DIN(N__47190),
            .DOUT(N__47189),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__47191),
            .PADOUT(N__47190),
            .PADIN(N__47189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__47182),
            .DIN(N__47181),
            .DOUT(N__47180),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__47182),
            .PADOUT(N__47181),
            .PADIN(N__47180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__47173),
            .DIN(N__47172),
            .DOUT(N__47171),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__47173),
            .PADOUT(N__47172),
            .PADIN(N__47171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21351),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__47164),
            .DIN(N__47163),
            .DOUT(N__47162),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__47164),
            .PADOUT(N__47163),
            .PADIN(N__47162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__47155),
            .DIN(N__47154),
            .DOUT(N__47153),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__47155),
            .PADOUT(N__47154),
            .PADIN(N__47153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36021),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_iopad (
            .OE(N__47146),
            .DIN(N__47145),
            .DOUT(N__47144),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_preio (
            .PADOEN(N__47146),
            .PADOUT(N__47145),
            .PADIN(N__47144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_iopad (
            .OE(N__47137),
            .DIN(N__47136),
            .DOUT(N__47135),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_preio (
            .PADOEN(N__47137),
            .PADOUT(N__47136),
            .PADIN(N__47135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__47128),
            .DIN(N__47127),
            .DOUT(N__47126),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__47128),
            .PADOUT(N__47127),
            .PADIN(N__47126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__47119),
            .DIN(N__47118),
            .DOUT(N__47117),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__47119),
            .PADOUT(N__47118),
            .PADIN(N__47117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33021),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__47110),
            .DIN(N__47109),
            .DOUT(N__47108),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__47110),
            .PADOUT(N__47109),
            .PADIN(N__47108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25611),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__47101),
            .DIN(N__47100),
            .DOUT(N__47099),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__47101),
            .PADOUT(N__47100),
            .PADIN(N__47099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__47092),
            .DIN(N__47091),
            .DOUT(N__47090),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__47092),
            .PADOUT(N__47091),
            .PADIN(N__47090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26148),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11252 (
            .O(N__47073),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__11251 (
            .O(N__47070),
            .I(N__47066));
    InMux I__11250 (
            .O(N__47069),
            .I(N__47063));
    LocalMux I__11249 (
            .O(N__47066),
            .I(N__47056));
    LocalMux I__11248 (
            .O(N__47063),
            .I(N__47053));
    InMux I__11247 (
            .O(N__47062),
            .I(N__47044));
    InMux I__11246 (
            .O(N__47061),
            .I(N__47044));
    InMux I__11245 (
            .O(N__47060),
            .I(N__47044));
    InMux I__11244 (
            .O(N__47059),
            .I(N__47044));
    Span4Mux_v I__11243 (
            .O(N__47056),
            .I(N__47041));
    Span12Mux_v I__11242 (
            .O(N__47053),
            .I(N__47038));
    LocalMux I__11241 (
            .O(N__47044),
            .I(N__47035));
    Odrv4 I__11240 (
            .O(N__47041),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__11239 (
            .O(N__47038),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__11238 (
            .O(N__47035),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__11237 (
            .O(N__47028),
            .I(N__47025));
    LocalMux I__11236 (
            .O(N__47025),
            .I(N__47022));
    Span4Mux_h I__11235 (
            .O(N__47022),
            .I(N__47017));
    InMux I__11234 (
            .O(N__47021),
            .I(N__47014));
    InMux I__11233 (
            .O(N__47020),
            .I(N__47011));
    Odrv4 I__11232 (
            .O(N__47017),
            .I(\phase_controller_inst1.stoper_hc.N_453 ));
    LocalMux I__11231 (
            .O(N__47014),
            .I(\phase_controller_inst1.stoper_hc.N_453 ));
    LocalMux I__11230 (
            .O(N__47011),
            .I(\phase_controller_inst1.stoper_hc.N_453 ));
    CascadeMux I__11229 (
            .O(N__47004),
            .I(N__47001));
    InMux I__11228 (
            .O(N__47001),
            .I(N__46998));
    LocalMux I__11227 (
            .O(N__46998),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__11226 (
            .O(N__46995),
            .I(N__46991));
    CascadeMux I__11225 (
            .O(N__46994),
            .I(N__46988));
    LocalMux I__11224 (
            .O(N__46991),
            .I(N__46985));
    InMux I__11223 (
            .O(N__46988),
            .I(N__46979));
    Span4Mux_h I__11222 (
            .O(N__46985),
            .I(N__46976));
    InMux I__11221 (
            .O(N__46984),
            .I(N__46973));
    InMux I__11220 (
            .O(N__46983),
            .I(N__46970));
    InMux I__11219 (
            .O(N__46982),
            .I(N__46967));
    LocalMux I__11218 (
            .O(N__46979),
            .I(measured_delay_hc_16));
    Odrv4 I__11217 (
            .O(N__46976),
            .I(measured_delay_hc_16));
    LocalMux I__11216 (
            .O(N__46973),
            .I(measured_delay_hc_16));
    LocalMux I__11215 (
            .O(N__46970),
            .I(measured_delay_hc_16));
    LocalMux I__11214 (
            .O(N__46967),
            .I(measured_delay_hc_16));
    CascadeMux I__11213 (
            .O(N__46956),
            .I(N__46953));
    InMux I__11212 (
            .O(N__46953),
            .I(N__46950));
    LocalMux I__11211 (
            .O(N__46950),
            .I(N__46947));
    Odrv4 I__11210 (
            .O(N__46947),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__11209 (
            .O(N__46944),
            .I(N__46931));
    CascadeMux I__11208 (
            .O(N__46943),
            .I(N__46928));
    CascadeMux I__11207 (
            .O(N__46942),
            .I(N__46925));
    CascadeMux I__11206 (
            .O(N__46941),
            .I(N__46922));
    InMux I__11205 (
            .O(N__46940),
            .I(N__46896));
    InMux I__11204 (
            .O(N__46939),
            .I(N__46896));
    InMux I__11203 (
            .O(N__46938),
            .I(N__46896));
    InMux I__11202 (
            .O(N__46937),
            .I(N__46896));
    InMux I__11201 (
            .O(N__46936),
            .I(N__46896));
    InMux I__11200 (
            .O(N__46935),
            .I(N__46896));
    InMux I__11199 (
            .O(N__46934),
            .I(N__46893));
    InMux I__11198 (
            .O(N__46931),
            .I(N__46873));
    InMux I__11197 (
            .O(N__46928),
            .I(N__46873));
    InMux I__11196 (
            .O(N__46925),
            .I(N__46873));
    InMux I__11195 (
            .O(N__46922),
            .I(N__46873));
    InMux I__11194 (
            .O(N__46921),
            .I(N__46873));
    InMux I__11193 (
            .O(N__46920),
            .I(N__46873));
    InMux I__11192 (
            .O(N__46919),
            .I(N__46873));
    InMux I__11191 (
            .O(N__46918),
            .I(N__46873));
    InMux I__11190 (
            .O(N__46917),
            .I(N__46868));
    InMux I__11189 (
            .O(N__46916),
            .I(N__46868));
    InMux I__11188 (
            .O(N__46915),
            .I(N__46853));
    InMux I__11187 (
            .O(N__46914),
            .I(N__46853));
    InMux I__11186 (
            .O(N__46913),
            .I(N__46853));
    InMux I__11185 (
            .O(N__46912),
            .I(N__46853));
    InMux I__11184 (
            .O(N__46911),
            .I(N__46853));
    InMux I__11183 (
            .O(N__46910),
            .I(N__46853));
    InMux I__11182 (
            .O(N__46909),
            .I(N__46853));
    LocalMux I__11181 (
            .O(N__46896),
            .I(N__46850));
    LocalMux I__11180 (
            .O(N__46893),
            .I(N__46847));
    InMux I__11179 (
            .O(N__46892),
            .I(N__46837));
    InMux I__11178 (
            .O(N__46891),
            .I(N__46837));
    InMux I__11177 (
            .O(N__46890),
            .I(N__46837));
    LocalMux I__11176 (
            .O(N__46873),
            .I(N__46825));
    LocalMux I__11175 (
            .O(N__46868),
            .I(N__46822));
    LocalMux I__11174 (
            .O(N__46853),
            .I(N__46815));
    Span4Mux_h I__11173 (
            .O(N__46850),
            .I(N__46815));
    Span4Mux_h I__11172 (
            .O(N__46847),
            .I(N__46815));
    InMux I__11171 (
            .O(N__46846),
            .I(N__46808));
    InMux I__11170 (
            .O(N__46845),
            .I(N__46808));
    InMux I__11169 (
            .O(N__46844),
            .I(N__46808));
    LocalMux I__11168 (
            .O(N__46837),
            .I(N__46805));
    InMux I__11167 (
            .O(N__46836),
            .I(N__46792));
    InMux I__11166 (
            .O(N__46835),
            .I(N__46792));
    InMux I__11165 (
            .O(N__46834),
            .I(N__46792));
    InMux I__11164 (
            .O(N__46833),
            .I(N__46792));
    InMux I__11163 (
            .O(N__46832),
            .I(N__46792));
    InMux I__11162 (
            .O(N__46831),
            .I(N__46792));
    InMux I__11161 (
            .O(N__46830),
            .I(N__46784));
    InMux I__11160 (
            .O(N__46829),
            .I(N__46784));
    InMux I__11159 (
            .O(N__46828),
            .I(N__46784));
    Span4Mux_v I__11158 (
            .O(N__46825),
            .I(N__46781));
    Span4Mux_h I__11157 (
            .O(N__46822),
            .I(N__46776));
    Span4Mux_v I__11156 (
            .O(N__46815),
            .I(N__46776));
    LocalMux I__11155 (
            .O(N__46808),
            .I(N__46769));
    Span4Mux_h I__11154 (
            .O(N__46805),
            .I(N__46769));
    LocalMux I__11153 (
            .O(N__46792),
            .I(N__46769));
    InMux I__11152 (
            .O(N__46791),
            .I(N__46766));
    LocalMux I__11151 (
            .O(N__46784),
            .I(\phase_controller_inst1.stoper_hc.N_449 ));
    Odrv4 I__11150 (
            .O(N__46781),
            .I(\phase_controller_inst1.stoper_hc.N_449 ));
    Odrv4 I__11149 (
            .O(N__46776),
            .I(\phase_controller_inst1.stoper_hc.N_449 ));
    Odrv4 I__11148 (
            .O(N__46769),
            .I(\phase_controller_inst1.stoper_hc.N_449 ));
    LocalMux I__11147 (
            .O(N__46766),
            .I(\phase_controller_inst1.stoper_hc.N_449 ));
    CascadeMux I__11146 (
            .O(N__46755),
            .I(N__46751));
    InMux I__11145 (
            .O(N__46754),
            .I(N__46748));
    InMux I__11144 (
            .O(N__46751),
            .I(N__46743));
    LocalMux I__11143 (
            .O(N__46748),
            .I(N__46740));
    InMux I__11142 (
            .O(N__46747),
            .I(N__46735));
    InMux I__11141 (
            .O(N__46746),
            .I(N__46735));
    LocalMux I__11140 (
            .O(N__46743),
            .I(N__46726));
    Span4Mux_v I__11139 (
            .O(N__46740),
            .I(N__46721));
    LocalMux I__11138 (
            .O(N__46735),
            .I(N__46721));
    CascadeMux I__11137 (
            .O(N__46734),
            .I(N__46718));
    InMux I__11136 (
            .O(N__46733),
            .I(N__46703));
    InMux I__11135 (
            .O(N__46732),
            .I(N__46703));
    InMux I__11134 (
            .O(N__46731),
            .I(N__46703));
    InMux I__11133 (
            .O(N__46730),
            .I(N__46703));
    InMux I__11132 (
            .O(N__46729),
            .I(N__46698));
    Span4Mux_v I__11131 (
            .O(N__46726),
            .I(N__46693));
    Span4Mux_h I__11130 (
            .O(N__46721),
            .I(N__46693));
    InMux I__11129 (
            .O(N__46718),
            .I(N__46686));
    InMux I__11128 (
            .O(N__46717),
            .I(N__46686));
    InMux I__11127 (
            .O(N__46716),
            .I(N__46686));
    InMux I__11126 (
            .O(N__46715),
            .I(N__46681));
    InMux I__11125 (
            .O(N__46714),
            .I(N__46681));
    InMux I__11124 (
            .O(N__46713),
            .I(N__46678));
    InMux I__11123 (
            .O(N__46712),
            .I(N__46675));
    LocalMux I__11122 (
            .O(N__46703),
            .I(N__46672));
    InMux I__11121 (
            .O(N__46702),
            .I(N__46667));
    InMux I__11120 (
            .O(N__46701),
            .I(N__46667));
    LocalMux I__11119 (
            .O(N__46698),
            .I(N__46664));
    Odrv4 I__11118 (
            .O(N__46693),
            .I(measured_delay_hc_31));
    LocalMux I__11117 (
            .O(N__46686),
            .I(measured_delay_hc_31));
    LocalMux I__11116 (
            .O(N__46681),
            .I(measured_delay_hc_31));
    LocalMux I__11115 (
            .O(N__46678),
            .I(measured_delay_hc_31));
    LocalMux I__11114 (
            .O(N__46675),
            .I(measured_delay_hc_31));
    Odrv4 I__11113 (
            .O(N__46672),
            .I(measured_delay_hc_31));
    LocalMux I__11112 (
            .O(N__46667),
            .I(measured_delay_hc_31));
    Odrv4 I__11111 (
            .O(N__46664),
            .I(measured_delay_hc_31));
    InMux I__11110 (
            .O(N__46647),
            .I(N__46644));
    LocalMux I__11109 (
            .O(N__46644),
            .I(N__46638));
    InMux I__11108 (
            .O(N__46643),
            .I(N__46634));
    InMux I__11107 (
            .O(N__46642),
            .I(N__46631));
    CascadeMux I__11106 (
            .O(N__46641),
            .I(N__46628));
    Span4Mux_h I__11105 (
            .O(N__46638),
            .I(N__46625));
    InMux I__11104 (
            .O(N__46637),
            .I(N__46622));
    LocalMux I__11103 (
            .O(N__46634),
            .I(N__46619));
    LocalMux I__11102 (
            .O(N__46631),
            .I(N__46616));
    InMux I__11101 (
            .O(N__46628),
            .I(N__46613));
    Span4Mux_v I__11100 (
            .O(N__46625),
            .I(N__46610));
    LocalMux I__11099 (
            .O(N__46622),
            .I(N__46607));
    Span4Mux_v I__11098 (
            .O(N__46619),
            .I(N__46602));
    Span4Mux_h I__11097 (
            .O(N__46616),
            .I(N__46602));
    LocalMux I__11096 (
            .O(N__46613),
            .I(measured_delay_hc_17));
    Odrv4 I__11095 (
            .O(N__46610),
            .I(measured_delay_hc_17));
    Odrv12 I__11094 (
            .O(N__46607),
            .I(measured_delay_hc_17));
    Odrv4 I__11093 (
            .O(N__46602),
            .I(measured_delay_hc_17));
    CascadeMux I__11092 (
            .O(N__46593),
            .I(N__46590));
    InMux I__11091 (
            .O(N__46590),
            .I(N__46587));
    LocalMux I__11090 (
            .O(N__46587),
            .I(N__46584));
    Odrv4 I__11089 (
            .O(N__46584),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    CEMux I__11088 (
            .O(N__46581),
            .I(N__46574));
    CEMux I__11087 (
            .O(N__46580),
            .I(N__46571));
    CEMux I__11086 (
            .O(N__46579),
            .I(N__46568));
    CEMux I__11085 (
            .O(N__46578),
            .I(N__46565));
    CEMux I__11084 (
            .O(N__46577),
            .I(N__46562));
    LocalMux I__11083 (
            .O(N__46574),
            .I(N__46558));
    LocalMux I__11082 (
            .O(N__46571),
            .I(N__46555));
    LocalMux I__11081 (
            .O(N__46568),
            .I(N__46552));
    LocalMux I__11080 (
            .O(N__46565),
            .I(N__46549));
    LocalMux I__11079 (
            .O(N__46562),
            .I(N__46546));
    CEMux I__11078 (
            .O(N__46561),
            .I(N__46543));
    Span4Mux_v I__11077 (
            .O(N__46558),
            .I(N__46540));
    Span4Mux_v I__11076 (
            .O(N__46555),
            .I(N__46535));
    Span4Mux_h I__11075 (
            .O(N__46552),
            .I(N__46535));
    Span4Mux_v I__11074 (
            .O(N__46549),
            .I(N__46528));
    Span4Mux_h I__11073 (
            .O(N__46546),
            .I(N__46528));
    LocalMux I__11072 (
            .O(N__46543),
            .I(N__46528));
    Span4Mux_h I__11071 (
            .O(N__46540),
            .I(N__46523));
    Span4Mux_h I__11070 (
            .O(N__46535),
            .I(N__46523));
    Span4Mux_v I__11069 (
            .O(N__46528),
            .I(N__46520));
    Odrv4 I__11068 (
            .O(N__46523),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__11067 (
            .O(N__46520),
            .I(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ));
    InMux I__11066 (
            .O(N__46515),
            .I(N__46511));
    InMux I__11065 (
            .O(N__46514),
            .I(N__46508));
    LocalMux I__11064 (
            .O(N__46511),
            .I(N__46505));
    LocalMux I__11063 (
            .O(N__46508),
            .I(measured_delay_hc_25));
    Odrv4 I__11062 (
            .O(N__46505),
            .I(measured_delay_hc_25));
    CascadeMux I__11061 (
            .O(N__46500),
            .I(N__46488));
    CascadeMux I__11060 (
            .O(N__46499),
            .I(N__46485));
    CascadeMux I__11059 (
            .O(N__46498),
            .I(N__46478));
    CascadeMux I__11058 (
            .O(N__46497),
            .I(N__46475));
    CascadeMux I__11057 (
            .O(N__46496),
            .I(N__46470));
    CascadeMux I__11056 (
            .O(N__46495),
            .I(N__46466));
    CascadeMux I__11055 (
            .O(N__46494),
            .I(N__46462));
    CascadeMux I__11054 (
            .O(N__46493),
            .I(N__46456));
    CascadeMux I__11053 (
            .O(N__46492),
            .I(N__46453));
    InMux I__11052 (
            .O(N__46491),
            .I(N__46440));
    InMux I__11051 (
            .O(N__46488),
            .I(N__46440));
    InMux I__11050 (
            .O(N__46485),
            .I(N__46440));
    InMux I__11049 (
            .O(N__46484),
            .I(N__46440));
    InMux I__11048 (
            .O(N__46483),
            .I(N__46434));
    InMux I__11047 (
            .O(N__46482),
            .I(N__46434));
    InMux I__11046 (
            .O(N__46481),
            .I(N__46423));
    InMux I__11045 (
            .O(N__46478),
            .I(N__46423));
    InMux I__11044 (
            .O(N__46475),
            .I(N__46423));
    InMux I__11043 (
            .O(N__46474),
            .I(N__46423));
    InMux I__11042 (
            .O(N__46473),
            .I(N__46423));
    InMux I__11041 (
            .O(N__46470),
            .I(N__46414));
    InMux I__11040 (
            .O(N__46469),
            .I(N__46414));
    InMux I__11039 (
            .O(N__46466),
            .I(N__46414));
    InMux I__11038 (
            .O(N__46465),
            .I(N__46414));
    InMux I__11037 (
            .O(N__46462),
            .I(N__46409));
    InMux I__11036 (
            .O(N__46461),
            .I(N__46409));
    InMux I__11035 (
            .O(N__46460),
            .I(N__46406));
    InMux I__11034 (
            .O(N__46459),
            .I(N__46395));
    InMux I__11033 (
            .O(N__46456),
            .I(N__46395));
    InMux I__11032 (
            .O(N__46453),
            .I(N__46395));
    InMux I__11031 (
            .O(N__46452),
            .I(N__46395));
    InMux I__11030 (
            .O(N__46451),
            .I(N__46395));
    CascadeMux I__11029 (
            .O(N__46450),
            .I(N__46392));
    CascadeMux I__11028 (
            .O(N__46449),
            .I(N__46389));
    LocalMux I__11027 (
            .O(N__46440),
            .I(N__46384));
    InMux I__11026 (
            .O(N__46439),
            .I(N__46381));
    LocalMux I__11025 (
            .O(N__46434),
            .I(N__46375));
    LocalMux I__11024 (
            .O(N__46423),
            .I(N__46370));
    LocalMux I__11023 (
            .O(N__46414),
            .I(N__46370));
    LocalMux I__11022 (
            .O(N__46409),
            .I(N__46367));
    LocalMux I__11021 (
            .O(N__46406),
            .I(N__46362));
    LocalMux I__11020 (
            .O(N__46395),
            .I(N__46362));
    InMux I__11019 (
            .O(N__46392),
            .I(N__46353));
    InMux I__11018 (
            .O(N__46389),
            .I(N__46353));
    InMux I__11017 (
            .O(N__46388),
            .I(N__46353));
    InMux I__11016 (
            .O(N__46387),
            .I(N__46353));
    Span4Mux_v I__11015 (
            .O(N__46384),
            .I(N__46347));
    LocalMux I__11014 (
            .O(N__46381),
            .I(N__46347));
    InMux I__11013 (
            .O(N__46380),
            .I(N__46340));
    InMux I__11012 (
            .O(N__46379),
            .I(N__46340));
    InMux I__11011 (
            .O(N__46378),
            .I(N__46340));
    Span4Mux_h I__11010 (
            .O(N__46375),
            .I(N__46335));
    Span4Mux_h I__11009 (
            .O(N__46370),
            .I(N__46335));
    Span4Mux_v I__11008 (
            .O(N__46367),
            .I(N__46328));
    Span4Mux_h I__11007 (
            .O(N__46362),
            .I(N__46328));
    LocalMux I__11006 (
            .O(N__46353),
            .I(N__46328));
    InMux I__11005 (
            .O(N__46352),
            .I(N__46325));
    Span4Mux_v I__11004 (
            .O(N__46347),
            .I(N__46320));
    LocalMux I__11003 (
            .O(N__46340),
            .I(N__46320));
    Odrv4 I__11002 (
            .O(N__46335),
            .I(\delay_measurement_inst.N_312 ));
    Odrv4 I__11001 (
            .O(N__46328),
            .I(\delay_measurement_inst.N_312 ));
    LocalMux I__11000 (
            .O(N__46325),
            .I(\delay_measurement_inst.N_312 ));
    Odrv4 I__10999 (
            .O(N__46320),
            .I(\delay_measurement_inst.N_312 ));
    CascadeMux I__10998 (
            .O(N__46311),
            .I(N__46308));
    InMux I__10997 (
            .O(N__46308),
            .I(N__46305));
    LocalMux I__10996 (
            .O(N__46305),
            .I(N__46301));
    InMux I__10995 (
            .O(N__46304),
            .I(N__46298));
    Span4Mux_v I__10994 (
            .O(N__46301),
            .I(N__46293));
    LocalMux I__10993 (
            .O(N__46298),
            .I(N__46293));
    Span4Mux_h I__10992 (
            .O(N__46293),
            .I(N__46289));
    InMux I__10991 (
            .O(N__46292),
            .I(N__46286));
    Odrv4 I__10990 (
            .O(N__46289),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    LocalMux I__10989 (
            .O(N__46286),
            .I(\delay_measurement_inst.elapsed_time_hc_2 ));
    InMux I__10988 (
            .O(N__46281),
            .I(N__46256));
    InMux I__10987 (
            .O(N__46280),
            .I(N__46256));
    InMux I__10986 (
            .O(N__46279),
            .I(N__46256));
    InMux I__10985 (
            .O(N__46278),
            .I(N__46256));
    InMux I__10984 (
            .O(N__46277),
            .I(N__46243));
    InMux I__10983 (
            .O(N__46276),
            .I(N__46243));
    InMux I__10982 (
            .O(N__46275),
            .I(N__46232));
    InMux I__10981 (
            .O(N__46274),
            .I(N__46232));
    InMux I__10980 (
            .O(N__46273),
            .I(N__46232));
    InMux I__10979 (
            .O(N__46272),
            .I(N__46232));
    InMux I__10978 (
            .O(N__46271),
            .I(N__46232));
    InMux I__10977 (
            .O(N__46270),
            .I(N__46223));
    InMux I__10976 (
            .O(N__46269),
            .I(N__46223));
    InMux I__10975 (
            .O(N__46268),
            .I(N__46223));
    InMux I__10974 (
            .O(N__46267),
            .I(N__46223));
    InMux I__10973 (
            .O(N__46266),
            .I(N__46215));
    InMux I__10972 (
            .O(N__46265),
            .I(N__46215));
    LocalMux I__10971 (
            .O(N__46256),
            .I(N__46212));
    InMux I__10970 (
            .O(N__46255),
            .I(N__46209));
    InMux I__10969 (
            .O(N__46254),
            .I(N__46206));
    InMux I__10968 (
            .O(N__46253),
            .I(N__46193));
    InMux I__10967 (
            .O(N__46252),
            .I(N__46193));
    InMux I__10966 (
            .O(N__46251),
            .I(N__46193));
    InMux I__10965 (
            .O(N__46250),
            .I(N__46193));
    InMux I__10964 (
            .O(N__46249),
            .I(N__46193));
    InMux I__10963 (
            .O(N__46248),
            .I(N__46193));
    LocalMux I__10962 (
            .O(N__46243),
            .I(N__46190));
    LocalMux I__10961 (
            .O(N__46232),
            .I(N__46185));
    LocalMux I__10960 (
            .O(N__46223),
            .I(N__46185));
    InMux I__10959 (
            .O(N__46222),
            .I(N__46178));
    InMux I__10958 (
            .O(N__46221),
            .I(N__46178));
    InMux I__10957 (
            .O(N__46220),
            .I(N__46178));
    LocalMux I__10956 (
            .O(N__46215),
            .I(N__46171));
    Span4Mux_v I__10955 (
            .O(N__46212),
            .I(N__46166));
    LocalMux I__10954 (
            .O(N__46209),
            .I(N__46166));
    LocalMux I__10953 (
            .O(N__46206),
            .I(N__46163));
    LocalMux I__10952 (
            .O(N__46193),
            .I(N__46160));
    Span4Mux_h I__10951 (
            .O(N__46190),
            .I(N__46153));
    Span4Mux_h I__10950 (
            .O(N__46185),
            .I(N__46153));
    LocalMux I__10949 (
            .O(N__46178),
            .I(N__46153));
    InMux I__10948 (
            .O(N__46177),
            .I(N__46144));
    InMux I__10947 (
            .O(N__46176),
            .I(N__46144));
    InMux I__10946 (
            .O(N__46175),
            .I(N__46144));
    InMux I__10945 (
            .O(N__46174),
            .I(N__46144));
    Odrv12 I__10944 (
            .O(N__46171),
            .I(\delay_measurement_inst.N_298 ));
    Odrv4 I__10943 (
            .O(N__46166),
            .I(\delay_measurement_inst.N_298 ));
    Odrv4 I__10942 (
            .O(N__46163),
            .I(\delay_measurement_inst.N_298 ));
    Odrv4 I__10941 (
            .O(N__46160),
            .I(\delay_measurement_inst.N_298 ));
    Odrv4 I__10940 (
            .O(N__46153),
            .I(\delay_measurement_inst.N_298 ));
    LocalMux I__10939 (
            .O(N__46144),
            .I(\delay_measurement_inst.N_298 ));
    InMux I__10938 (
            .O(N__46131),
            .I(N__46125));
    InMux I__10937 (
            .O(N__46130),
            .I(N__46122));
    InMux I__10936 (
            .O(N__46129),
            .I(N__46119));
    InMux I__10935 (
            .O(N__46128),
            .I(N__46116));
    LocalMux I__10934 (
            .O(N__46125),
            .I(N__46113));
    LocalMux I__10933 (
            .O(N__46122),
            .I(N__46109));
    LocalMux I__10932 (
            .O(N__46119),
            .I(N__46106));
    LocalMux I__10931 (
            .O(N__46116),
            .I(N__46103));
    Span4Mux_h I__10930 (
            .O(N__46113),
            .I(N__46100));
    InMux I__10929 (
            .O(N__46112),
            .I(N__46097));
    Span4Mux_v I__10928 (
            .O(N__46109),
            .I(N__46094));
    Span4Mux_h I__10927 (
            .O(N__46106),
            .I(N__46091));
    Span4Mux_v I__10926 (
            .O(N__46103),
            .I(N__46086));
    Span4Mux_v I__10925 (
            .O(N__46100),
            .I(N__46086));
    LocalMux I__10924 (
            .O(N__46097),
            .I(measured_delay_hc_2));
    Odrv4 I__10923 (
            .O(N__46094),
            .I(measured_delay_hc_2));
    Odrv4 I__10922 (
            .O(N__46091),
            .I(measured_delay_hc_2));
    Odrv4 I__10921 (
            .O(N__46086),
            .I(measured_delay_hc_2));
    ClkMux I__10920 (
            .O(N__46077),
            .I(N__45627));
    ClkMux I__10919 (
            .O(N__46076),
            .I(N__45627));
    ClkMux I__10918 (
            .O(N__46075),
            .I(N__45627));
    ClkMux I__10917 (
            .O(N__46074),
            .I(N__45627));
    ClkMux I__10916 (
            .O(N__46073),
            .I(N__45627));
    ClkMux I__10915 (
            .O(N__46072),
            .I(N__45627));
    ClkMux I__10914 (
            .O(N__46071),
            .I(N__45627));
    ClkMux I__10913 (
            .O(N__46070),
            .I(N__45627));
    ClkMux I__10912 (
            .O(N__46069),
            .I(N__45627));
    ClkMux I__10911 (
            .O(N__46068),
            .I(N__45627));
    ClkMux I__10910 (
            .O(N__46067),
            .I(N__45627));
    ClkMux I__10909 (
            .O(N__46066),
            .I(N__45627));
    ClkMux I__10908 (
            .O(N__46065),
            .I(N__45627));
    ClkMux I__10907 (
            .O(N__46064),
            .I(N__45627));
    ClkMux I__10906 (
            .O(N__46063),
            .I(N__45627));
    ClkMux I__10905 (
            .O(N__46062),
            .I(N__45627));
    ClkMux I__10904 (
            .O(N__46061),
            .I(N__45627));
    ClkMux I__10903 (
            .O(N__46060),
            .I(N__45627));
    ClkMux I__10902 (
            .O(N__46059),
            .I(N__45627));
    ClkMux I__10901 (
            .O(N__46058),
            .I(N__45627));
    ClkMux I__10900 (
            .O(N__46057),
            .I(N__45627));
    ClkMux I__10899 (
            .O(N__46056),
            .I(N__45627));
    ClkMux I__10898 (
            .O(N__46055),
            .I(N__45627));
    ClkMux I__10897 (
            .O(N__46054),
            .I(N__45627));
    ClkMux I__10896 (
            .O(N__46053),
            .I(N__45627));
    ClkMux I__10895 (
            .O(N__46052),
            .I(N__45627));
    ClkMux I__10894 (
            .O(N__46051),
            .I(N__45627));
    ClkMux I__10893 (
            .O(N__46050),
            .I(N__45627));
    ClkMux I__10892 (
            .O(N__46049),
            .I(N__45627));
    ClkMux I__10891 (
            .O(N__46048),
            .I(N__45627));
    ClkMux I__10890 (
            .O(N__46047),
            .I(N__45627));
    ClkMux I__10889 (
            .O(N__46046),
            .I(N__45627));
    ClkMux I__10888 (
            .O(N__46045),
            .I(N__45627));
    ClkMux I__10887 (
            .O(N__46044),
            .I(N__45627));
    ClkMux I__10886 (
            .O(N__46043),
            .I(N__45627));
    ClkMux I__10885 (
            .O(N__46042),
            .I(N__45627));
    ClkMux I__10884 (
            .O(N__46041),
            .I(N__45627));
    ClkMux I__10883 (
            .O(N__46040),
            .I(N__45627));
    ClkMux I__10882 (
            .O(N__46039),
            .I(N__45627));
    ClkMux I__10881 (
            .O(N__46038),
            .I(N__45627));
    ClkMux I__10880 (
            .O(N__46037),
            .I(N__45627));
    ClkMux I__10879 (
            .O(N__46036),
            .I(N__45627));
    ClkMux I__10878 (
            .O(N__46035),
            .I(N__45627));
    ClkMux I__10877 (
            .O(N__46034),
            .I(N__45627));
    ClkMux I__10876 (
            .O(N__46033),
            .I(N__45627));
    ClkMux I__10875 (
            .O(N__46032),
            .I(N__45627));
    ClkMux I__10874 (
            .O(N__46031),
            .I(N__45627));
    ClkMux I__10873 (
            .O(N__46030),
            .I(N__45627));
    ClkMux I__10872 (
            .O(N__46029),
            .I(N__45627));
    ClkMux I__10871 (
            .O(N__46028),
            .I(N__45627));
    ClkMux I__10870 (
            .O(N__46027),
            .I(N__45627));
    ClkMux I__10869 (
            .O(N__46026),
            .I(N__45627));
    ClkMux I__10868 (
            .O(N__46025),
            .I(N__45627));
    ClkMux I__10867 (
            .O(N__46024),
            .I(N__45627));
    ClkMux I__10866 (
            .O(N__46023),
            .I(N__45627));
    ClkMux I__10865 (
            .O(N__46022),
            .I(N__45627));
    ClkMux I__10864 (
            .O(N__46021),
            .I(N__45627));
    ClkMux I__10863 (
            .O(N__46020),
            .I(N__45627));
    ClkMux I__10862 (
            .O(N__46019),
            .I(N__45627));
    ClkMux I__10861 (
            .O(N__46018),
            .I(N__45627));
    ClkMux I__10860 (
            .O(N__46017),
            .I(N__45627));
    ClkMux I__10859 (
            .O(N__46016),
            .I(N__45627));
    ClkMux I__10858 (
            .O(N__46015),
            .I(N__45627));
    ClkMux I__10857 (
            .O(N__46014),
            .I(N__45627));
    ClkMux I__10856 (
            .O(N__46013),
            .I(N__45627));
    ClkMux I__10855 (
            .O(N__46012),
            .I(N__45627));
    ClkMux I__10854 (
            .O(N__46011),
            .I(N__45627));
    ClkMux I__10853 (
            .O(N__46010),
            .I(N__45627));
    ClkMux I__10852 (
            .O(N__46009),
            .I(N__45627));
    ClkMux I__10851 (
            .O(N__46008),
            .I(N__45627));
    ClkMux I__10850 (
            .O(N__46007),
            .I(N__45627));
    ClkMux I__10849 (
            .O(N__46006),
            .I(N__45627));
    ClkMux I__10848 (
            .O(N__46005),
            .I(N__45627));
    ClkMux I__10847 (
            .O(N__46004),
            .I(N__45627));
    ClkMux I__10846 (
            .O(N__46003),
            .I(N__45627));
    ClkMux I__10845 (
            .O(N__46002),
            .I(N__45627));
    ClkMux I__10844 (
            .O(N__46001),
            .I(N__45627));
    ClkMux I__10843 (
            .O(N__46000),
            .I(N__45627));
    ClkMux I__10842 (
            .O(N__45999),
            .I(N__45627));
    ClkMux I__10841 (
            .O(N__45998),
            .I(N__45627));
    ClkMux I__10840 (
            .O(N__45997),
            .I(N__45627));
    ClkMux I__10839 (
            .O(N__45996),
            .I(N__45627));
    ClkMux I__10838 (
            .O(N__45995),
            .I(N__45627));
    ClkMux I__10837 (
            .O(N__45994),
            .I(N__45627));
    ClkMux I__10836 (
            .O(N__45993),
            .I(N__45627));
    ClkMux I__10835 (
            .O(N__45992),
            .I(N__45627));
    ClkMux I__10834 (
            .O(N__45991),
            .I(N__45627));
    ClkMux I__10833 (
            .O(N__45990),
            .I(N__45627));
    ClkMux I__10832 (
            .O(N__45989),
            .I(N__45627));
    ClkMux I__10831 (
            .O(N__45988),
            .I(N__45627));
    ClkMux I__10830 (
            .O(N__45987),
            .I(N__45627));
    ClkMux I__10829 (
            .O(N__45986),
            .I(N__45627));
    ClkMux I__10828 (
            .O(N__45985),
            .I(N__45627));
    ClkMux I__10827 (
            .O(N__45984),
            .I(N__45627));
    ClkMux I__10826 (
            .O(N__45983),
            .I(N__45627));
    ClkMux I__10825 (
            .O(N__45982),
            .I(N__45627));
    ClkMux I__10824 (
            .O(N__45981),
            .I(N__45627));
    ClkMux I__10823 (
            .O(N__45980),
            .I(N__45627));
    ClkMux I__10822 (
            .O(N__45979),
            .I(N__45627));
    ClkMux I__10821 (
            .O(N__45978),
            .I(N__45627));
    ClkMux I__10820 (
            .O(N__45977),
            .I(N__45627));
    ClkMux I__10819 (
            .O(N__45976),
            .I(N__45627));
    ClkMux I__10818 (
            .O(N__45975),
            .I(N__45627));
    ClkMux I__10817 (
            .O(N__45974),
            .I(N__45627));
    ClkMux I__10816 (
            .O(N__45973),
            .I(N__45627));
    ClkMux I__10815 (
            .O(N__45972),
            .I(N__45627));
    ClkMux I__10814 (
            .O(N__45971),
            .I(N__45627));
    ClkMux I__10813 (
            .O(N__45970),
            .I(N__45627));
    ClkMux I__10812 (
            .O(N__45969),
            .I(N__45627));
    ClkMux I__10811 (
            .O(N__45968),
            .I(N__45627));
    ClkMux I__10810 (
            .O(N__45967),
            .I(N__45627));
    ClkMux I__10809 (
            .O(N__45966),
            .I(N__45627));
    ClkMux I__10808 (
            .O(N__45965),
            .I(N__45627));
    ClkMux I__10807 (
            .O(N__45964),
            .I(N__45627));
    ClkMux I__10806 (
            .O(N__45963),
            .I(N__45627));
    ClkMux I__10805 (
            .O(N__45962),
            .I(N__45627));
    ClkMux I__10804 (
            .O(N__45961),
            .I(N__45627));
    ClkMux I__10803 (
            .O(N__45960),
            .I(N__45627));
    ClkMux I__10802 (
            .O(N__45959),
            .I(N__45627));
    ClkMux I__10801 (
            .O(N__45958),
            .I(N__45627));
    ClkMux I__10800 (
            .O(N__45957),
            .I(N__45627));
    ClkMux I__10799 (
            .O(N__45956),
            .I(N__45627));
    ClkMux I__10798 (
            .O(N__45955),
            .I(N__45627));
    ClkMux I__10797 (
            .O(N__45954),
            .I(N__45627));
    ClkMux I__10796 (
            .O(N__45953),
            .I(N__45627));
    ClkMux I__10795 (
            .O(N__45952),
            .I(N__45627));
    ClkMux I__10794 (
            .O(N__45951),
            .I(N__45627));
    ClkMux I__10793 (
            .O(N__45950),
            .I(N__45627));
    ClkMux I__10792 (
            .O(N__45949),
            .I(N__45627));
    ClkMux I__10791 (
            .O(N__45948),
            .I(N__45627));
    ClkMux I__10790 (
            .O(N__45947),
            .I(N__45627));
    ClkMux I__10789 (
            .O(N__45946),
            .I(N__45627));
    ClkMux I__10788 (
            .O(N__45945),
            .I(N__45627));
    ClkMux I__10787 (
            .O(N__45944),
            .I(N__45627));
    ClkMux I__10786 (
            .O(N__45943),
            .I(N__45627));
    ClkMux I__10785 (
            .O(N__45942),
            .I(N__45627));
    ClkMux I__10784 (
            .O(N__45941),
            .I(N__45627));
    ClkMux I__10783 (
            .O(N__45940),
            .I(N__45627));
    ClkMux I__10782 (
            .O(N__45939),
            .I(N__45627));
    ClkMux I__10781 (
            .O(N__45938),
            .I(N__45627));
    ClkMux I__10780 (
            .O(N__45937),
            .I(N__45627));
    ClkMux I__10779 (
            .O(N__45936),
            .I(N__45627));
    ClkMux I__10778 (
            .O(N__45935),
            .I(N__45627));
    ClkMux I__10777 (
            .O(N__45934),
            .I(N__45627));
    ClkMux I__10776 (
            .O(N__45933),
            .I(N__45627));
    ClkMux I__10775 (
            .O(N__45932),
            .I(N__45627));
    ClkMux I__10774 (
            .O(N__45931),
            .I(N__45627));
    ClkMux I__10773 (
            .O(N__45930),
            .I(N__45627));
    ClkMux I__10772 (
            .O(N__45929),
            .I(N__45627));
    ClkMux I__10771 (
            .O(N__45928),
            .I(N__45627));
    GlobalMux I__10770 (
            .O(N__45627),
            .I(clk_100mhz_0));
    CascadeMux I__10769 (
            .O(N__45624),
            .I(N__45615));
    CascadeMux I__10768 (
            .O(N__45623),
            .I(N__45612));
    InMux I__10767 (
            .O(N__45622),
            .I(N__45609));
    InMux I__10766 (
            .O(N__45621),
            .I(N__45606));
    InMux I__10765 (
            .O(N__45620),
            .I(N__45603));
    InMux I__10764 (
            .O(N__45619),
            .I(N__45600));
    InMux I__10763 (
            .O(N__45618),
            .I(N__45597));
    InMux I__10762 (
            .O(N__45615),
            .I(N__45594));
    InMux I__10761 (
            .O(N__45612),
            .I(N__45591));
    LocalMux I__10760 (
            .O(N__45609),
            .I(N__45588));
    LocalMux I__10759 (
            .O(N__45606),
            .I(N__45585));
    LocalMux I__10758 (
            .O(N__45603),
            .I(N__45582));
    LocalMux I__10757 (
            .O(N__45600),
            .I(N__45536));
    LocalMux I__10756 (
            .O(N__45597),
            .I(N__45470));
    LocalMux I__10755 (
            .O(N__45594),
            .I(N__45462));
    LocalMux I__10754 (
            .O(N__45591),
            .I(N__45449));
    Glb2LocalMux I__10753 (
            .O(N__45588),
            .I(N__45165));
    Glb2LocalMux I__10752 (
            .O(N__45585),
            .I(N__45165));
    Glb2LocalMux I__10751 (
            .O(N__45582),
            .I(N__45165));
    SRMux I__10750 (
            .O(N__45581),
            .I(N__45165));
    SRMux I__10749 (
            .O(N__45580),
            .I(N__45165));
    SRMux I__10748 (
            .O(N__45579),
            .I(N__45165));
    SRMux I__10747 (
            .O(N__45578),
            .I(N__45165));
    SRMux I__10746 (
            .O(N__45577),
            .I(N__45165));
    SRMux I__10745 (
            .O(N__45576),
            .I(N__45165));
    SRMux I__10744 (
            .O(N__45575),
            .I(N__45165));
    SRMux I__10743 (
            .O(N__45574),
            .I(N__45165));
    SRMux I__10742 (
            .O(N__45573),
            .I(N__45165));
    SRMux I__10741 (
            .O(N__45572),
            .I(N__45165));
    SRMux I__10740 (
            .O(N__45571),
            .I(N__45165));
    SRMux I__10739 (
            .O(N__45570),
            .I(N__45165));
    SRMux I__10738 (
            .O(N__45569),
            .I(N__45165));
    SRMux I__10737 (
            .O(N__45568),
            .I(N__45165));
    SRMux I__10736 (
            .O(N__45567),
            .I(N__45165));
    SRMux I__10735 (
            .O(N__45566),
            .I(N__45165));
    SRMux I__10734 (
            .O(N__45565),
            .I(N__45165));
    SRMux I__10733 (
            .O(N__45564),
            .I(N__45165));
    SRMux I__10732 (
            .O(N__45563),
            .I(N__45165));
    SRMux I__10731 (
            .O(N__45562),
            .I(N__45165));
    SRMux I__10730 (
            .O(N__45561),
            .I(N__45165));
    SRMux I__10729 (
            .O(N__45560),
            .I(N__45165));
    SRMux I__10728 (
            .O(N__45559),
            .I(N__45165));
    SRMux I__10727 (
            .O(N__45558),
            .I(N__45165));
    SRMux I__10726 (
            .O(N__45557),
            .I(N__45165));
    SRMux I__10725 (
            .O(N__45556),
            .I(N__45165));
    SRMux I__10724 (
            .O(N__45555),
            .I(N__45165));
    SRMux I__10723 (
            .O(N__45554),
            .I(N__45165));
    SRMux I__10722 (
            .O(N__45553),
            .I(N__45165));
    SRMux I__10721 (
            .O(N__45552),
            .I(N__45165));
    SRMux I__10720 (
            .O(N__45551),
            .I(N__45165));
    SRMux I__10719 (
            .O(N__45550),
            .I(N__45165));
    SRMux I__10718 (
            .O(N__45549),
            .I(N__45165));
    SRMux I__10717 (
            .O(N__45548),
            .I(N__45165));
    SRMux I__10716 (
            .O(N__45547),
            .I(N__45165));
    SRMux I__10715 (
            .O(N__45546),
            .I(N__45165));
    SRMux I__10714 (
            .O(N__45545),
            .I(N__45165));
    SRMux I__10713 (
            .O(N__45544),
            .I(N__45165));
    SRMux I__10712 (
            .O(N__45543),
            .I(N__45165));
    SRMux I__10711 (
            .O(N__45542),
            .I(N__45165));
    SRMux I__10710 (
            .O(N__45541),
            .I(N__45165));
    SRMux I__10709 (
            .O(N__45540),
            .I(N__45165));
    SRMux I__10708 (
            .O(N__45539),
            .I(N__45165));
    Glb2LocalMux I__10707 (
            .O(N__45536),
            .I(N__45165));
    SRMux I__10706 (
            .O(N__45535),
            .I(N__45165));
    SRMux I__10705 (
            .O(N__45534),
            .I(N__45165));
    SRMux I__10704 (
            .O(N__45533),
            .I(N__45165));
    SRMux I__10703 (
            .O(N__45532),
            .I(N__45165));
    SRMux I__10702 (
            .O(N__45531),
            .I(N__45165));
    SRMux I__10701 (
            .O(N__45530),
            .I(N__45165));
    SRMux I__10700 (
            .O(N__45529),
            .I(N__45165));
    SRMux I__10699 (
            .O(N__45528),
            .I(N__45165));
    SRMux I__10698 (
            .O(N__45527),
            .I(N__45165));
    SRMux I__10697 (
            .O(N__45526),
            .I(N__45165));
    SRMux I__10696 (
            .O(N__45525),
            .I(N__45165));
    SRMux I__10695 (
            .O(N__45524),
            .I(N__45165));
    SRMux I__10694 (
            .O(N__45523),
            .I(N__45165));
    SRMux I__10693 (
            .O(N__45522),
            .I(N__45165));
    SRMux I__10692 (
            .O(N__45521),
            .I(N__45165));
    SRMux I__10691 (
            .O(N__45520),
            .I(N__45165));
    SRMux I__10690 (
            .O(N__45519),
            .I(N__45165));
    SRMux I__10689 (
            .O(N__45518),
            .I(N__45165));
    SRMux I__10688 (
            .O(N__45517),
            .I(N__45165));
    SRMux I__10687 (
            .O(N__45516),
            .I(N__45165));
    SRMux I__10686 (
            .O(N__45515),
            .I(N__45165));
    SRMux I__10685 (
            .O(N__45514),
            .I(N__45165));
    SRMux I__10684 (
            .O(N__45513),
            .I(N__45165));
    SRMux I__10683 (
            .O(N__45512),
            .I(N__45165));
    SRMux I__10682 (
            .O(N__45511),
            .I(N__45165));
    SRMux I__10681 (
            .O(N__45510),
            .I(N__45165));
    SRMux I__10680 (
            .O(N__45509),
            .I(N__45165));
    SRMux I__10679 (
            .O(N__45508),
            .I(N__45165));
    SRMux I__10678 (
            .O(N__45507),
            .I(N__45165));
    SRMux I__10677 (
            .O(N__45506),
            .I(N__45165));
    SRMux I__10676 (
            .O(N__45505),
            .I(N__45165));
    SRMux I__10675 (
            .O(N__45504),
            .I(N__45165));
    SRMux I__10674 (
            .O(N__45503),
            .I(N__45165));
    SRMux I__10673 (
            .O(N__45502),
            .I(N__45165));
    SRMux I__10672 (
            .O(N__45501),
            .I(N__45165));
    SRMux I__10671 (
            .O(N__45500),
            .I(N__45165));
    SRMux I__10670 (
            .O(N__45499),
            .I(N__45165));
    SRMux I__10669 (
            .O(N__45498),
            .I(N__45165));
    SRMux I__10668 (
            .O(N__45497),
            .I(N__45165));
    SRMux I__10667 (
            .O(N__45496),
            .I(N__45165));
    SRMux I__10666 (
            .O(N__45495),
            .I(N__45165));
    SRMux I__10665 (
            .O(N__45494),
            .I(N__45165));
    SRMux I__10664 (
            .O(N__45493),
            .I(N__45165));
    SRMux I__10663 (
            .O(N__45492),
            .I(N__45165));
    SRMux I__10662 (
            .O(N__45491),
            .I(N__45165));
    SRMux I__10661 (
            .O(N__45490),
            .I(N__45165));
    SRMux I__10660 (
            .O(N__45489),
            .I(N__45165));
    SRMux I__10659 (
            .O(N__45488),
            .I(N__45165));
    SRMux I__10658 (
            .O(N__45487),
            .I(N__45165));
    SRMux I__10657 (
            .O(N__45486),
            .I(N__45165));
    SRMux I__10656 (
            .O(N__45485),
            .I(N__45165));
    SRMux I__10655 (
            .O(N__45484),
            .I(N__45165));
    SRMux I__10654 (
            .O(N__45483),
            .I(N__45165));
    SRMux I__10653 (
            .O(N__45482),
            .I(N__45165));
    SRMux I__10652 (
            .O(N__45481),
            .I(N__45165));
    SRMux I__10651 (
            .O(N__45480),
            .I(N__45165));
    SRMux I__10650 (
            .O(N__45479),
            .I(N__45165));
    SRMux I__10649 (
            .O(N__45478),
            .I(N__45165));
    SRMux I__10648 (
            .O(N__45477),
            .I(N__45165));
    SRMux I__10647 (
            .O(N__45476),
            .I(N__45165));
    SRMux I__10646 (
            .O(N__45475),
            .I(N__45165));
    SRMux I__10645 (
            .O(N__45474),
            .I(N__45165));
    SRMux I__10644 (
            .O(N__45473),
            .I(N__45165));
    Glb2LocalMux I__10643 (
            .O(N__45470),
            .I(N__45165));
    SRMux I__10642 (
            .O(N__45469),
            .I(N__45165));
    SRMux I__10641 (
            .O(N__45468),
            .I(N__45165));
    SRMux I__10640 (
            .O(N__45467),
            .I(N__45165));
    SRMux I__10639 (
            .O(N__45466),
            .I(N__45165));
    SRMux I__10638 (
            .O(N__45465),
            .I(N__45165));
    Glb2LocalMux I__10637 (
            .O(N__45462),
            .I(N__45165));
    SRMux I__10636 (
            .O(N__45461),
            .I(N__45165));
    SRMux I__10635 (
            .O(N__45460),
            .I(N__45165));
    SRMux I__10634 (
            .O(N__45459),
            .I(N__45165));
    SRMux I__10633 (
            .O(N__45458),
            .I(N__45165));
    SRMux I__10632 (
            .O(N__45457),
            .I(N__45165));
    SRMux I__10631 (
            .O(N__45456),
            .I(N__45165));
    SRMux I__10630 (
            .O(N__45455),
            .I(N__45165));
    SRMux I__10629 (
            .O(N__45454),
            .I(N__45165));
    SRMux I__10628 (
            .O(N__45453),
            .I(N__45165));
    SRMux I__10627 (
            .O(N__45452),
            .I(N__45165));
    Glb2LocalMux I__10626 (
            .O(N__45449),
            .I(N__45165));
    SRMux I__10625 (
            .O(N__45448),
            .I(N__45165));
    SRMux I__10624 (
            .O(N__45447),
            .I(N__45165));
    SRMux I__10623 (
            .O(N__45446),
            .I(N__45165));
    SRMux I__10622 (
            .O(N__45445),
            .I(N__45165));
    SRMux I__10621 (
            .O(N__45444),
            .I(N__45165));
    SRMux I__10620 (
            .O(N__45443),
            .I(N__45165));
    SRMux I__10619 (
            .O(N__45442),
            .I(N__45165));
    SRMux I__10618 (
            .O(N__45441),
            .I(N__45165));
    SRMux I__10617 (
            .O(N__45440),
            .I(N__45165));
    GlobalMux I__10616 (
            .O(N__45165),
            .I(N__45162));
    gio2CtrlBuf I__10615 (
            .O(N__45162),
            .I(red_c_g));
    CascadeMux I__10614 (
            .O(N__45159),
            .I(N__45156));
    InMux I__10613 (
            .O(N__45156),
            .I(N__45153));
    LocalMux I__10612 (
            .O(N__45153),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__10611 (
            .O(N__45150),
            .I(N__45146));
    InMux I__10610 (
            .O(N__45149),
            .I(N__45143));
    LocalMux I__10609 (
            .O(N__45146),
            .I(N__45140));
    LocalMux I__10608 (
            .O(N__45143),
            .I(N__45137));
    Odrv4 I__10607 (
            .O(N__45140),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__10606 (
            .O(N__45137),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__10605 (
            .O(N__45132),
            .I(N__45129));
    LocalMux I__10604 (
            .O(N__45129),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__10603 (
            .O(N__45126),
            .I(N__45123));
    LocalMux I__10602 (
            .O(N__45123),
            .I(N__45119));
    InMux I__10601 (
            .O(N__45122),
            .I(N__45116));
    Span4Mux_v I__10600 (
            .O(N__45119),
            .I(N__45111));
    LocalMux I__10599 (
            .O(N__45116),
            .I(N__45111));
    Odrv4 I__10598 (
            .O(N__45111),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__10597 (
            .O(N__45108),
            .I(N__45105));
    InMux I__10596 (
            .O(N__45105),
            .I(N__45102));
    LocalMux I__10595 (
            .O(N__45102),
            .I(N__45099));
    Odrv4 I__10594 (
            .O(N__45099),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__10593 (
            .O(N__45096),
            .I(N__45093));
    LocalMux I__10592 (
            .O(N__45093),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__10591 (
            .O(N__45090),
            .I(N__45087));
    LocalMux I__10590 (
            .O(N__45087),
            .I(N__45084));
    Span4Mux_h I__10589 (
            .O(N__45084),
            .I(N__45081));
    Odrv4 I__10588 (
            .O(N__45081),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__10587 (
            .O(N__45078),
            .I(N__45074));
    InMux I__10586 (
            .O(N__45077),
            .I(N__45071));
    LocalMux I__10585 (
            .O(N__45074),
            .I(N__45068));
    LocalMux I__10584 (
            .O(N__45071),
            .I(N__45065));
    Span4Mux_v I__10583 (
            .O(N__45068),
            .I(N__45062));
    Odrv4 I__10582 (
            .O(N__45065),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__10581 (
            .O(N__45062),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__10580 (
            .O(N__45057),
            .I(N__45054));
    InMux I__10579 (
            .O(N__45054),
            .I(N__45051));
    LocalMux I__10578 (
            .O(N__45051),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__10577 (
            .O(N__45048),
            .I(N__45045));
    InMux I__10576 (
            .O(N__45045),
            .I(N__45042));
    LocalMux I__10575 (
            .O(N__45042),
            .I(N__45039));
    Odrv4 I__10574 (
            .O(N__45039),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__10573 (
            .O(N__45036),
            .I(N__45033));
    LocalMux I__10572 (
            .O(N__45033),
            .I(N__45029));
    InMux I__10571 (
            .O(N__45032),
            .I(N__45026));
    Span4Mux_h I__10570 (
            .O(N__45029),
            .I(N__45023));
    LocalMux I__10569 (
            .O(N__45026),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__10568 (
            .O(N__45023),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__10567 (
            .O(N__45018),
            .I(N__45015));
    LocalMux I__10566 (
            .O(N__45015),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__10565 (
            .O(N__45012),
            .I(N__45009));
    LocalMux I__10564 (
            .O(N__45009),
            .I(N__45005));
    InMux I__10563 (
            .O(N__45008),
            .I(N__45002));
    Span4Mux_v I__10562 (
            .O(N__45005),
            .I(N__44999));
    LocalMux I__10561 (
            .O(N__45002),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__10560 (
            .O(N__44999),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__10559 (
            .O(N__44994),
            .I(N__44991));
    LocalMux I__10558 (
            .O(N__44991),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ));
    InMux I__10557 (
            .O(N__44988),
            .I(N__44984));
    InMux I__10556 (
            .O(N__44987),
            .I(N__44981));
    LocalMux I__10555 (
            .O(N__44984),
            .I(N__44978));
    LocalMux I__10554 (
            .O(N__44981),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__10553 (
            .O(N__44978),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__10552 (
            .O(N__44973),
            .I(N__44970));
    LocalMux I__10551 (
            .O(N__44970),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ));
    CascadeMux I__10550 (
            .O(N__44967),
            .I(N__44964));
    InMux I__10549 (
            .O(N__44964),
            .I(N__44961));
    LocalMux I__10548 (
            .O(N__44961),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__10547 (
            .O(N__44958),
            .I(N__44954));
    InMux I__10546 (
            .O(N__44957),
            .I(N__44951));
    LocalMux I__10545 (
            .O(N__44954),
            .I(N__44948));
    LocalMux I__10544 (
            .O(N__44951),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__10543 (
            .O(N__44948),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__10542 (
            .O(N__44943),
            .I(N__44940));
    LocalMux I__10541 (
            .O(N__44940),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ));
    InMux I__10540 (
            .O(N__44937),
            .I(N__44933));
    InMux I__10539 (
            .O(N__44936),
            .I(N__44930));
    LocalMux I__10538 (
            .O(N__44933),
            .I(N__44927));
    LocalMux I__10537 (
            .O(N__44930),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__10536 (
            .O(N__44927),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__10535 (
            .O(N__44922),
            .I(N__44919));
    LocalMux I__10534 (
            .O(N__44919),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ));
    CascadeMux I__10533 (
            .O(N__44916),
            .I(N__44913));
    InMux I__10532 (
            .O(N__44913),
            .I(N__44910));
    LocalMux I__10531 (
            .O(N__44910),
            .I(N__44907));
    Odrv4 I__10530 (
            .O(N__44907),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    InMux I__10529 (
            .O(N__44904),
            .I(N__44901));
    LocalMux I__10528 (
            .O(N__44901),
            .I(N__44897));
    InMux I__10527 (
            .O(N__44900),
            .I(N__44894));
    Odrv4 I__10526 (
            .O(N__44897),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__10525 (
            .O(N__44894),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__10524 (
            .O(N__44889),
            .I(N__44886));
    LocalMux I__10523 (
            .O(N__44886),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__10522 (
            .O(N__44883),
            .I(N__44880));
    LocalMux I__10521 (
            .O(N__44880),
            .I(N__44876));
    InMux I__10520 (
            .O(N__44879),
            .I(N__44873));
    Odrv4 I__10519 (
            .O(N__44876),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__10518 (
            .O(N__44873),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__10517 (
            .O(N__44868),
            .I(N__44865));
    InMux I__10516 (
            .O(N__44865),
            .I(N__44862));
    LocalMux I__10515 (
            .O(N__44862),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    InMux I__10514 (
            .O(N__44859),
            .I(N__44856));
    LocalMux I__10513 (
            .O(N__44856),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__10512 (
            .O(N__44853),
            .I(N__44850));
    LocalMux I__10511 (
            .O(N__44850),
            .I(N__44846));
    InMux I__10510 (
            .O(N__44849),
            .I(N__44843));
    Odrv4 I__10509 (
            .O(N__44846),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__10508 (
            .O(N__44843),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__10507 (
            .O(N__44838),
            .I(N__44835));
    InMux I__10506 (
            .O(N__44835),
            .I(N__44832));
    LocalMux I__10505 (
            .O(N__44832),
            .I(N__44829));
    Odrv4 I__10504 (
            .O(N__44829),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__10503 (
            .O(N__44826),
            .I(N__44823));
    LocalMux I__10502 (
            .O(N__44823),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__10501 (
            .O(N__44820),
            .I(N__44817));
    LocalMux I__10500 (
            .O(N__44817),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    InMux I__10499 (
            .O(N__44814),
            .I(N__44810));
    InMux I__10498 (
            .O(N__44813),
            .I(N__44807));
    LocalMux I__10497 (
            .O(N__44810),
            .I(N__44804));
    LocalMux I__10496 (
            .O(N__44807),
            .I(N__44801));
    Odrv12 I__10495 (
            .O(N__44804),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__10494 (
            .O(N__44801),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__10493 (
            .O(N__44796),
            .I(N__44793));
    InMux I__10492 (
            .O(N__44793),
            .I(N__44790));
    LocalMux I__10491 (
            .O(N__44790),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__10490 (
            .O(N__44787),
            .I(N__44784));
    InMux I__10489 (
            .O(N__44784),
            .I(N__44781));
    LocalMux I__10488 (
            .O(N__44781),
            .I(N__44778));
    Odrv4 I__10487 (
            .O(N__44778),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__10486 (
            .O(N__44775),
            .I(N__44771));
    InMux I__10485 (
            .O(N__44774),
            .I(N__44768));
    LocalMux I__10484 (
            .O(N__44771),
            .I(N__44765));
    LocalMux I__10483 (
            .O(N__44768),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__10482 (
            .O(N__44765),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__10481 (
            .O(N__44760),
            .I(N__44757));
    LocalMux I__10480 (
            .O(N__44757),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__10479 (
            .O(N__44754),
            .I(N__44751));
    InMux I__10478 (
            .O(N__44751),
            .I(N__44748));
    LocalMux I__10477 (
            .O(N__44748),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__10476 (
            .O(N__44745),
            .I(N__44741));
    InMux I__10475 (
            .O(N__44744),
            .I(N__44738));
    LocalMux I__10474 (
            .O(N__44741),
            .I(N__44735));
    LocalMux I__10473 (
            .O(N__44738),
            .I(N__44730));
    Span12Mux_v I__10472 (
            .O(N__44735),
            .I(N__44730));
    Odrv12 I__10471 (
            .O(N__44730),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__10470 (
            .O(N__44727),
            .I(N__44724));
    LocalMux I__10469 (
            .O(N__44724),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__10468 (
            .O(N__44721),
            .I(N__44718));
    InMux I__10467 (
            .O(N__44718),
            .I(N__44715));
    LocalMux I__10466 (
            .O(N__44715),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__10465 (
            .O(N__44712),
            .I(N__44709));
    LocalMux I__10464 (
            .O(N__44709),
            .I(N__44705));
    InMux I__10463 (
            .O(N__44708),
            .I(N__44702));
    Span4Mux_v I__10462 (
            .O(N__44705),
            .I(N__44699));
    LocalMux I__10461 (
            .O(N__44702),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__10460 (
            .O(N__44699),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__10459 (
            .O(N__44694),
            .I(N__44691));
    LocalMux I__10458 (
            .O(N__44691),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__10457 (
            .O(N__44688),
            .I(N__44685));
    InMux I__10456 (
            .O(N__44685),
            .I(N__44682));
    LocalMux I__10455 (
            .O(N__44682),
            .I(N__44679));
    Odrv12 I__10454 (
            .O(N__44679),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ));
    InMux I__10453 (
            .O(N__44676),
            .I(N__44673));
    LocalMux I__10452 (
            .O(N__44673),
            .I(N__44670));
    Odrv4 I__10451 (
            .O(N__44670),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ));
    InMux I__10450 (
            .O(N__44667),
            .I(N__44657));
    InMux I__10449 (
            .O(N__44666),
            .I(N__44657));
    CascadeMux I__10448 (
            .O(N__44665),
            .I(N__44654));
    CascadeMux I__10447 (
            .O(N__44664),
            .I(N__44650));
    CascadeMux I__10446 (
            .O(N__44663),
            .I(N__44636));
    CascadeMux I__10445 (
            .O(N__44662),
            .I(N__44633));
    LocalMux I__10444 (
            .O(N__44657),
            .I(N__44628));
    InMux I__10443 (
            .O(N__44654),
            .I(N__44623));
    InMux I__10442 (
            .O(N__44653),
            .I(N__44623));
    InMux I__10441 (
            .O(N__44650),
            .I(N__44606));
    InMux I__10440 (
            .O(N__44649),
            .I(N__44606));
    InMux I__10439 (
            .O(N__44648),
            .I(N__44606));
    InMux I__10438 (
            .O(N__44647),
            .I(N__44606));
    InMux I__10437 (
            .O(N__44646),
            .I(N__44606));
    InMux I__10436 (
            .O(N__44645),
            .I(N__44606));
    InMux I__10435 (
            .O(N__44644),
            .I(N__44606));
    InMux I__10434 (
            .O(N__44643),
            .I(N__44606));
    CascadeMux I__10433 (
            .O(N__44642),
            .I(N__44603));
    CascadeMux I__10432 (
            .O(N__44641),
            .I(N__44600));
    CascadeMux I__10431 (
            .O(N__44640),
            .I(N__44597));
    InMux I__10430 (
            .O(N__44639),
            .I(N__44586));
    InMux I__10429 (
            .O(N__44636),
            .I(N__44586));
    InMux I__10428 (
            .O(N__44633),
            .I(N__44586));
    InMux I__10427 (
            .O(N__44632),
            .I(N__44586));
    InMux I__10426 (
            .O(N__44631),
            .I(N__44586));
    Span4Mux_h I__10425 (
            .O(N__44628),
            .I(N__44579));
    LocalMux I__10424 (
            .O(N__44623),
            .I(N__44579));
    LocalMux I__10423 (
            .O(N__44606),
            .I(N__44576));
    InMux I__10422 (
            .O(N__44603),
            .I(N__44569));
    InMux I__10421 (
            .O(N__44600),
            .I(N__44569));
    InMux I__10420 (
            .O(N__44597),
            .I(N__44569));
    LocalMux I__10419 (
            .O(N__44586),
            .I(N__44566));
    InMux I__10418 (
            .O(N__44585),
            .I(N__44561));
    InMux I__10417 (
            .O(N__44584),
            .I(N__44561));
    Span4Mux_v I__10416 (
            .O(N__44579),
            .I(N__44554));
    Span4Mux_v I__10415 (
            .O(N__44576),
            .I(N__44554));
    LocalMux I__10414 (
            .O(N__44569),
            .I(N__44547));
    Span4Mux_v I__10413 (
            .O(N__44566),
            .I(N__44547));
    LocalMux I__10412 (
            .O(N__44561),
            .I(N__44547));
    InMux I__10411 (
            .O(N__44560),
            .I(N__44544));
    CascadeMux I__10410 (
            .O(N__44559),
            .I(N__44541));
    Span4Mux_h I__10409 (
            .O(N__44554),
            .I(N__44538));
    Span4Mux_v I__10408 (
            .O(N__44547),
            .I(N__44535));
    LocalMux I__10407 (
            .O(N__44544),
            .I(N__44532));
    InMux I__10406 (
            .O(N__44541),
            .I(N__44529));
    Span4Mux_v I__10405 (
            .O(N__44538),
            .I(N__44526));
    Span4Mux_v I__10404 (
            .O(N__44535),
            .I(N__44523));
    Span12Mux_h I__10403 (
            .O(N__44532),
            .I(N__44520));
    LocalMux I__10402 (
            .O(N__44529),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__10401 (
            .O(N__44526),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__10400 (
            .O(N__44523),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv12 I__10399 (
            .O(N__44520),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    CascadeMux I__10398 (
            .O(N__44511),
            .I(N__44502));
    CascadeMux I__10397 (
            .O(N__44510),
            .I(N__44499));
    CascadeMux I__10396 (
            .O(N__44509),
            .I(N__44496));
    CascadeMux I__10395 (
            .O(N__44508),
            .I(N__44493));
    CascadeMux I__10394 (
            .O(N__44507),
            .I(N__44486));
    CascadeMux I__10393 (
            .O(N__44506),
            .I(N__44483));
    CascadeMux I__10392 (
            .O(N__44505),
            .I(N__44478));
    InMux I__10391 (
            .O(N__44502),
            .I(N__44455));
    InMux I__10390 (
            .O(N__44499),
            .I(N__44455));
    InMux I__10389 (
            .O(N__44496),
            .I(N__44455));
    InMux I__10388 (
            .O(N__44493),
            .I(N__44455));
    InMux I__10387 (
            .O(N__44492),
            .I(N__44455));
    InMux I__10386 (
            .O(N__44491),
            .I(N__44455));
    InMux I__10385 (
            .O(N__44490),
            .I(N__44455));
    InMux I__10384 (
            .O(N__44489),
            .I(N__44455));
    InMux I__10383 (
            .O(N__44486),
            .I(N__44446));
    InMux I__10382 (
            .O(N__44483),
            .I(N__44446));
    InMux I__10381 (
            .O(N__44482),
            .I(N__44446));
    InMux I__10380 (
            .O(N__44481),
            .I(N__44446));
    InMux I__10379 (
            .O(N__44478),
            .I(N__44441));
    InMux I__10378 (
            .O(N__44477),
            .I(N__44434));
    InMux I__10377 (
            .O(N__44476),
            .I(N__44434));
    InMux I__10376 (
            .O(N__44475),
            .I(N__44434));
    CascadeMux I__10375 (
            .O(N__44474),
            .I(N__44430));
    InMux I__10374 (
            .O(N__44473),
            .I(N__44423));
    InMux I__10373 (
            .O(N__44472),
            .I(N__44423));
    LocalMux I__10372 (
            .O(N__44455),
            .I(N__44418));
    LocalMux I__10371 (
            .O(N__44446),
            .I(N__44418));
    InMux I__10370 (
            .O(N__44445),
            .I(N__44413));
    InMux I__10369 (
            .O(N__44444),
            .I(N__44413));
    LocalMux I__10368 (
            .O(N__44441),
            .I(N__44410));
    LocalMux I__10367 (
            .O(N__44434),
            .I(N__44407));
    InMux I__10366 (
            .O(N__44433),
            .I(N__44404));
    InMux I__10365 (
            .O(N__44430),
            .I(N__44397));
    InMux I__10364 (
            .O(N__44429),
            .I(N__44397));
    InMux I__10363 (
            .O(N__44428),
            .I(N__44397));
    LocalMux I__10362 (
            .O(N__44423),
            .I(N__44394));
    Span4Mux_v I__10361 (
            .O(N__44418),
            .I(N__44391));
    LocalMux I__10360 (
            .O(N__44413),
            .I(N__44380));
    Span4Mux_v I__10359 (
            .O(N__44410),
            .I(N__44380));
    Span4Mux_h I__10358 (
            .O(N__44407),
            .I(N__44380));
    LocalMux I__10357 (
            .O(N__44404),
            .I(N__44380));
    LocalMux I__10356 (
            .O(N__44397),
            .I(N__44380));
    Odrv4 I__10355 (
            .O(N__44394),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__10354 (
            .O(N__44391),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__10353 (
            .O(N__44380),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__10352 (
            .O(N__44373),
            .I(N__44370));
    InMux I__10351 (
            .O(N__44370),
            .I(N__44367));
    LocalMux I__10350 (
            .O(N__44367),
            .I(N__44364));
    Span4Mux_v I__10349 (
            .O(N__44364),
            .I(N__44361));
    Odrv4 I__10348 (
            .O(N__44361),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ));
    CascadeMux I__10347 (
            .O(N__44358),
            .I(N__44354));
    InMux I__10346 (
            .O(N__44357),
            .I(N__44334));
    InMux I__10345 (
            .O(N__44354),
            .I(N__44331));
    InMux I__10344 (
            .O(N__44353),
            .I(N__44314));
    InMux I__10343 (
            .O(N__44352),
            .I(N__44314));
    InMux I__10342 (
            .O(N__44351),
            .I(N__44314));
    InMux I__10341 (
            .O(N__44350),
            .I(N__44314));
    InMux I__10340 (
            .O(N__44349),
            .I(N__44314));
    InMux I__10339 (
            .O(N__44348),
            .I(N__44314));
    InMux I__10338 (
            .O(N__44347),
            .I(N__44314));
    InMux I__10337 (
            .O(N__44346),
            .I(N__44314));
    InMux I__10336 (
            .O(N__44345),
            .I(N__44303));
    InMux I__10335 (
            .O(N__44344),
            .I(N__44303));
    InMux I__10334 (
            .O(N__44343),
            .I(N__44303));
    InMux I__10333 (
            .O(N__44342),
            .I(N__44303));
    InMux I__10332 (
            .O(N__44341),
            .I(N__44303));
    CascadeMux I__10331 (
            .O(N__44340),
            .I(N__44295));
    InMux I__10330 (
            .O(N__44339),
            .I(N__44288));
    InMux I__10329 (
            .O(N__44338),
            .I(N__44288));
    InMux I__10328 (
            .O(N__44337),
            .I(N__44288));
    LocalMux I__10327 (
            .O(N__44334),
            .I(N__44283));
    LocalMux I__10326 (
            .O(N__44331),
            .I(N__44283));
    LocalMux I__10325 (
            .O(N__44314),
            .I(N__44278));
    LocalMux I__10324 (
            .O(N__44303),
            .I(N__44278));
    InMux I__10323 (
            .O(N__44302),
            .I(N__44275));
    InMux I__10322 (
            .O(N__44301),
            .I(N__44268));
    InMux I__10321 (
            .O(N__44300),
            .I(N__44268));
    InMux I__10320 (
            .O(N__44299),
            .I(N__44268));
    InMux I__10319 (
            .O(N__44298),
            .I(N__44263));
    InMux I__10318 (
            .O(N__44295),
            .I(N__44263));
    LocalMux I__10317 (
            .O(N__44288),
            .I(N__44252));
    Span4Mux_v I__10316 (
            .O(N__44283),
            .I(N__44252));
    Span4Mux_v I__10315 (
            .O(N__44278),
            .I(N__44252));
    LocalMux I__10314 (
            .O(N__44275),
            .I(N__44252));
    LocalMux I__10313 (
            .O(N__44268),
            .I(N__44252));
    LocalMux I__10312 (
            .O(N__44263),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10311 (
            .O(N__44252),
            .I(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__10310 (
            .O(N__44247),
            .I(N__44244));
    InMux I__10309 (
            .O(N__44244),
            .I(N__44241));
    LocalMux I__10308 (
            .O(N__44241),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__10307 (
            .O(N__44238),
            .I(N__44235));
    InMux I__10306 (
            .O(N__44235),
            .I(N__44232));
    LocalMux I__10305 (
            .O(N__44232),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__10304 (
            .O(N__44229),
            .I(N__44225));
    InMux I__10303 (
            .O(N__44228),
            .I(N__44222));
    InMux I__10302 (
            .O(N__44225),
            .I(N__44218));
    LocalMux I__10301 (
            .O(N__44222),
            .I(N__44215));
    InMux I__10300 (
            .O(N__44221),
            .I(N__44212));
    LocalMux I__10299 (
            .O(N__44218),
            .I(N__44207));
    Span12Mux_v I__10298 (
            .O(N__44215),
            .I(N__44207));
    LocalMux I__10297 (
            .O(N__44212),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv12 I__10296 (
            .O(N__44207),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__10295 (
            .O(N__44202),
            .I(N__44199));
    LocalMux I__10294 (
            .O(N__44199),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    CascadeMux I__10293 (
            .O(N__44196),
            .I(N__44193));
    InMux I__10292 (
            .O(N__44193),
            .I(N__44190));
    LocalMux I__10291 (
            .O(N__44190),
            .I(N__44187));
    Odrv4 I__10290 (
            .O(N__44187),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__10289 (
            .O(N__44184),
            .I(N__44181));
    LocalMux I__10288 (
            .O(N__44181),
            .I(N__44177));
    InMux I__10287 (
            .O(N__44180),
            .I(N__44174));
    Odrv12 I__10286 (
            .O(N__44177),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__10285 (
            .O(N__44174),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__10284 (
            .O(N__44169),
            .I(N__44166));
    LocalMux I__10283 (
            .O(N__44166),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__10282 (
            .O(N__44163),
            .I(N__44160));
    InMux I__10281 (
            .O(N__44160),
            .I(N__44157));
    LocalMux I__10280 (
            .O(N__44157),
            .I(N__44153));
    InMux I__10279 (
            .O(N__44156),
            .I(N__44150));
    Odrv4 I__10278 (
            .O(N__44153),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__10277 (
            .O(N__44150),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__10276 (
            .O(N__44145),
            .I(N__44142));
    InMux I__10275 (
            .O(N__44142),
            .I(N__44139));
    LocalMux I__10274 (
            .O(N__44139),
            .I(N__44136));
    Span4Mux_h I__10273 (
            .O(N__44136),
            .I(N__44133));
    Odrv4 I__10272 (
            .O(N__44133),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    InMux I__10271 (
            .O(N__44130),
            .I(N__44127));
    LocalMux I__10270 (
            .O(N__44127),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__10269 (
            .O(N__44124),
            .I(N__44121));
    InMux I__10268 (
            .O(N__44121),
            .I(N__44118));
    LocalMux I__10267 (
            .O(N__44118),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    InMux I__10266 (
            .O(N__44115),
            .I(N__44112));
    LocalMux I__10265 (
            .O(N__44112),
            .I(N__44108));
    InMux I__10264 (
            .O(N__44111),
            .I(N__44105));
    Odrv12 I__10263 (
            .O(N__44108),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__10262 (
            .O(N__44105),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__10261 (
            .O(N__44100),
            .I(N__44097));
    LocalMux I__10260 (
            .O(N__44097),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__10259 (
            .O(N__44094),
            .I(N__44091));
    LocalMux I__10258 (
            .O(N__44091),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ));
    InMux I__10257 (
            .O(N__44088),
            .I(bfn_18_15_0_));
    InMux I__10256 (
            .O(N__44085),
            .I(N__44082));
    LocalMux I__10255 (
            .O(N__44082),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ));
    InMux I__10254 (
            .O(N__44079),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__10253 (
            .O(N__44076),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__10252 (
            .O(N__44073),
            .I(N__44070));
    LocalMux I__10251 (
            .O(N__44070),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ));
    InMux I__10250 (
            .O(N__44067),
            .I(N__44064));
    LocalMux I__10249 (
            .O(N__44064),
            .I(N__44061));
    Odrv4 I__10248 (
            .O(N__44061),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ));
    CascadeMux I__10247 (
            .O(N__44058),
            .I(N__44055));
    InMux I__10246 (
            .O(N__44055),
            .I(N__44052));
    LocalMux I__10245 (
            .O(N__44052),
            .I(N__44049));
    Odrv4 I__10244 (
            .O(N__44049),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ));
    InMux I__10243 (
            .O(N__44046),
            .I(N__44043));
    LocalMux I__10242 (
            .O(N__44043),
            .I(N__44040));
    Odrv4 I__10241 (
            .O(N__44040),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ));
    InMux I__10240 (
            .O(N__44037),
            .I(N__44034));
    LocalMux I__10239 (
            .O(N__44034),
            .I(N__44031));
    Odrv4 I__10238 (
            .O(N__44031),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ));
    InMux I__10237 (
            .O(N__44028),
            .I(N__44025));
    LocalMux I__10236 (
            .O(N__44025),
            .I(N__44022));
    Odrv4 I__10235 (
            .O(N__44022),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ));
    InMux I__10234 (
            .O(N__44019),
            .I(N__44016));
    LocalMux I__10233 (
            .O(N__44016),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ));
    InMux I__10232 (
            .O(N__44013),
            .I(bfn_18_14_0_));
    InMux I__10231 (
            .O(N__44010),
            .I(N__44007));
    LocalMux I__10230 (
            .O(N__44007),
            .I(N__44004));
    Odrv12 I__10229 (
            .O(N__44004),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ));
    InMux I__10228 (
            .O(N__44001),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__10227 (
            .O(N__43998),
            .I(N__43995));
    LocalMux I__10226 (
            .O(N__43995),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ));
    InMux I__10225 (
            .O(N__43992),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__10224 (
            .O(N__43989),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__10223 (
            .O(N__43986),
            .I(N__43983));
    LocalMux I__10222 (
            .O(N__43983),
            .I(N__43980));
    Odrv4 I__10221 (
            .O(N__43980),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ));
    InMux I__10220 (
            .O(N__43977),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ));
    InMux I__10219 (
            .O(N__43974),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__10218 (
            .O(N__43971),
            .I(N__43968));
    LocalMux I__10217 (
            .O(N__43968),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ));
    InMux I__10216 (
            .O(N__43965),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__10215 (
            .O(N__43962),
            .I(N__43959));
    LocalMux I__10214 (
            .O(N__43959),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ));
    InMux I__10213 (
            .O(N__43956),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__10212 (
            .O(N__43953),
            .I(N__43949));
    CascadeMux I__10211 (
            .O(N__43952),
            .I(N__43946));
    LocalMux I__10210 (
            .O(N__43949),
            .I(N__43941));
    InMux I__10209 (
            .O(N__43946),
            .I(N__43936));
    InMux I__10208 (
            .O(N__43945),
            .I(N__43936));
    InMux I__10207 (
            .O(N__43944),
            .I(N__43933));
    Span4Mux_v I__10206 (
            .O(N__43941),
            .I(N__43928));
    LocalMux I__10205 (
            .O(N__43936),
            .I(N__43928));
    LocalMux I__10204 (
            .O(N__43933),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    Odrv4 I__10203 (
            .O(N__43928),
            .I(\phase_controller_inst2.stoper_hc.time_passed11 ));
    InMux I__10202 (
            .O(N__43923),
            .I(N__43920));
    LocalMux I__10201 (
            .O(N__43920),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ));
    InMux I__10200 (
            .O(N__43917),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__10199 (
            .O(N__43914),
            .I(N__43911));
    LocalMux I__10198 (
            .O(N__43911),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ));
    InMux I__10197 (
            .O(N__43908),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__10196 (
            .O(N__43905),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__10195 (
            .O(N__43902),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__10194 (
            .O(N__43899),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__10193 (
            .O(N__43896),
            .I(N__43893));
    LocalMux I__10192 (
            .O(N__43893),
            .I(N__43890));
    Odrv4 I__10191 (
            .O(N__43890),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ));
    InMux I__10190 (
            .O(N__43887),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__10189 (
            .O(N__43884),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__10188 (
            .O(N__43881),
            .I(N__43877));
    InMux I__10187 (
            .O(N__43880),
            .I(N__43874));
    LocalMux I__10186 (
            .O(N__43877),
            .I(N__43871));
    LocalMux I__10185 (
            .O(N__43874),
            .I(N__43867));
    Span4Mux_v I__10184 (
            .O(N__43871),
            .I(N__43864));
    InMux I__10183 (
            .O(N__43870),
            .I(N__43861));
    Odrv4 I__10182 (
            .O(N__43867),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__10181 (
            .O(N__43864),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__10180 (
            .O(N__43861),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__10179 (
            .O(N__43854),
            .I(N__43851));
    LocalMux I__10178 (
            .O(N__43851),
            .I(N__43847));
    CascadeMux I__10177 (
            .O(N__43850),
            .I(N__43844));
    Span4Mux_v I__10176 (
            .O(N__43847),
            .I(N__43841));
    InMux I__10175 (
            .O(N__43844),
            .I(N__43838));
    Span4Mux_v I__10174 (
            .O(N__43841),
            .I(N__43833));
    LocalMux I__10173 (
            .O(N__43838),
            .I(N__43833));
    Odrv4 I__10172 (
            .O(N__43833),
            .I(\delay_measurement_inst.elapsed_time_tr_1 ));
    CEMux I__10171 (
            .O(N__43830),
            .I(N__43812));
    CEMux I__10170 (
            .O(N__43829),
            .I(N__43812));
    CEMux I__10169 (
            .O(N__43828),
            .I(N__43812));
    CEMux I__10168 (
            .O(N__43827),
            .I(N__43812));
    CEMux I__10167 (
            .O(N__43826),
            .I(N__43812));
    CEMux I__10166 (
            .O(N__43825),
            .I(N__43812));
    GlobalMux I__10165 (
            .O(N__43812),
            .I(N__43809));
    gio2CtrlBuf I__10164 (
            .O(N__43809),
            .I(\delay_measurement_inst.delay_tr_timer.N_463_i_g ));
    CascadeMux I__10163 (
            .O(N__43806),
            .I(N__43802));
    InMux I__10162 (
            .O(N__43805),
            .I(N__43798));
    InMux I__10161 (
            .O(N__43802),
            .I(N__43793));
    InMux I__10160 (
            .O(N__43801),
            .I(N__43793));
    LocalMux I__10159 (
            .O(N__43798),
            .I(N__43790));
    LocalMux I__10158 (
            .O(N__43793),
            .I(N__43787));
    Span4Mux_h I__10157 (
            .O(N__43790),
            .I(N__43784));
    Span4Mux_h I__10156 (
            .O(N__43787),
            .I(N__43781));
    Odrv4 I__10155 (
            .O(N__43784),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    Odrv4 I__10154 (
            .O(N__43781),
            .I(\delay_measurement_inst.elapsed_time_tr_17 ));
    InMux I__10153 (
            .O(N__43776),
            .I(N__43772));
    InMux I__10152 (
            .O(N__43775),
            .I(N__43769));
    LocalMux I__10151 (
            .O(N__43772),
            .I(N__43766));
    LocalMux I__10150 (
            .O(N__43769),
            .I(N__43763));
    Span4Mux_v I__10149 (
            .O(N__43766),
            .I(N__43758));
    Span4Mux_v I__10148 (
            .O(N__43763),
            .I(N__43755));
    InMux I__10147 (
            .O(N__43762),
            .I(N__43750));
    InMux I__10146 (
            .O(N__43761),
            .I(N__43750));
    Span4Mux_h I__10145 (
            .O(N__43758),
            .I(N__43747));
    Span4Mux_h I__10144 (
            .O(N__43755),
            .I(N__43742));
    LocalMux I__10143 (
            .O(N__43750),
            .I(N__43742));
    Sp12to4 I__10142 (
            .O(N__43747),
            .I(N__43739));
    Span4Mux_h I__10141 (
            .O(N__43742),
            .I(N__43736));
    Odrv12 I__10140 (
            .O(N__43739),
            .I(measured_delay_tr_17));
    Odrv4 I__10139 (
            .O(N__43736),
            .I(measured_delay_tr_17));
    InMux I__10138 (
            .O(N__43731),
            .I(N__43723));
    InMux I__10137 (
            .O(N__43730),
            .I(N__43723));
    InMux I__10136 (
            .O(N__43729),
            .I(N__43716));
    InMux I__10135 (
            .O(N__43728),
            .I(N__43716));
    LocalMux I__10134 (
            .O(N__43723),
            .I(N__43713));
    InMux I__10133 (
            .O(N__43722),
            .I(N__43708));
    InMux I__10132 (
            .O(N__43721),
            .I(N__43708));
    LocalMux I__10131 (
            .O(N__43716),
            .I(N__43702));
    Span4Mux_h I__10130 (
            .O(N__43713),
            .I(N__43699));
    LocalMux I__10129 (
            .O(N__43708),
            .I(N__43696));
    InMux I__10128 (
            .O(N__43707),
            .I(N__43691));
    InMux I__10127 (
            .O(N__43706),
            .I(N__43691));
    InMux I__10126 (
            .O(N__43705),
            .I(N__43688));
    Odrv4 I__10125 (
            .O(N__43702),
            .I(\delay_measurement_inst.N_498 ));
    Odrv4 I__10124 (
            .O(N__43699),
            .I(\delay_measurement_inst.N_498 ));
    Odrv4 I__10123 (
            .O(N__43696),
            .I(\delay_measurement_inst.N_498 ));
    LocalMux I__10122 (
            .O(N__43691),
            .I(\delay_measurement_inst.N_498 ));
    LocalMux I__10121 (
            .O(N__43688),
            .I(\delay_measurement_inst.N_498 ));
    CascadeMux I__10120 (
            .O(N__43677),
            .I(N__43667));
    CascadeMux I__10119 (
            .O(N__43676),
            .I(N__43662));
    CascadeMux I__10118 (
            .O(N__43675),
            .I(N__43657));
    CascadeMux I__10117 (
            .O(N__43674),
            .I(N__43654));
    InMux I__10116 (
            .O(N__43673),
            .I(N__43649));
    InMux I__10115 (
            .O(N__43672),
            .I(N__43649));
    InMux I__10114 (
            .O(N__43671),
            .I(N__43636));
    InMux I__10113 (
            .O(N__43670),
            .I(N__43636));
    InMux I__10112 (
            .O(N__43667),
            .I(N__43636));
    InMux I__10111 (
            .O(N__43666),
            .I(N__43636));
    InMux I__10110 (
            .O(N__43665),
            .I(N__43636));
    InMux I__10109 (
            .O(N__43662),
            .I(N__43629));
    InMux I__10108 (
            .O(N__43661),
            .I(N__43629));
    InMux I__10107 (
            .O(N__43660),
            .I(N__43629));
    InMux I__10106 (
            .O(N__43657),
            .I(N__43626));
    InMux I__10105 (
            .O(N__43654),
            .I(N__43623));
    LocalMux I__10104 (
            .O(N__43649),
            .I(N__43620));
    InMux I__10103 (
            .O(N__43648),
            .I(N__43615));
    InMux I__10102 (
            .O(N__43647),
            .I(N__43615));
    LocalMux I__10101 (
            .O(N__43636),
            .I(N__43610));
    LocalMux I__10100 (
            .O(N__43629),
            .I(N__43610));
    LocalMux I__10099 (
            .O(N__43626),
            .I(N__43607));
    LocalMux I__10098 (
            .O(N__43623),
            .I(N__43604));
    Span4Mux_v I__10097 (
            .O(N__43620),
            .I(N__43601));
    LocalMux I__10096 (
            .O(N__43615),
            .I(N__43598));
    Span4Mux_h I__10095 (
            .O(N__43610),
            .I(N__43595));
    Span4Mux_v I__10094 (
            .O(N__43607),
            .I(N__43590));
    Span4Mux_v I__10093 (
            .O(N__43604),
            .I(N__43590));
    Odrv4 I__10092 (
            .O(N__43601),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv12 I__10091 (
            .O(N__43598),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__10090 (
            .O(N__43595),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__10089 (
            .O(N__43590),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    InMux I__10088 (
            .O(N__43581),
            .I(N__43578));
    LocalMux I__10087 (
            .O(N__43578),
            .I(N__43573));
    InMux I__10086 (
            .O(N__43577),
            .I(N__43568));
    InMux I__10085 (
            .O(N__43576),
            .I(N__43568));
    Span4Mux_h I__10084 (
            .O(N__43573),
            .I(N__43565));
    LocalMux I__10083 (
            .O(N__43568),
            .I(N__43562));
    Odrv4 I__10082 (
            .O(N__43565),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    Odrv4 I__10081 (
            .O(N__43562),
            .I(\delay_measurement_inst.elapsed_time_tr_18 ));
    InMux I__10080 (
            .O(N__43557),
            .I(N__43553));
    InMux I__10079 (
            .O(N__43556),
            .I(N__43550));
    LocalMux I__10078 (
            .O(N__43553),
            .I(N__43547));
    LocalMux I__10077 (
            .O(N__43550),
            .I(N__43544));
    Span4Mux_v I__10076 (
            .O(N__43547),
            .I(N__43539));
    Span4Mux_v I__10075 (
            .O(N__43544),
            .I(N__43536));
    InMux I__10074 (
            .O(N__43543),
            .I(N__43531));
    InMux I__10073 (
            .O(N__43542),
            .I(N__43531));
    Sp12to4 I__10072 (
            .O(N__43539),
            .I(N__43524));
    Sp12to4 I__10071 (
            .O(N__43536),
            .I(N__43524));
    LocalMux I__10070 (
            .O(N__43531),
            .I(N__43524));
    Odrv12 I__10069 (
            .O(N__43524),
            .I(measured_delay_tr_18));
    CEMux I__10068 (
            .O(N__43521),
            .I(N__43516));
    CEMux I__10067 (
            .O(N__43520),
            .I(N__43512));
    CEMux I__10066 (
            .O(N__43519),
            .I(N__43508));
    LocalMux I__10065 (
            .O(N__43516),
            .I(N__43505));
    CEMux I__10064 (
            .O(N__43515),
            .I(N__43502));
    LocalMux I__10063 (
            .O(N__43512),
            .I(N__43499));
    CEMux I__10062 (
            .O(N__43511),
            .I(N__43496));
    LocalMux I__10061 (
            .O(N__43508),
            .I(N__43493));
    Span4Mux_h I__10060 (
            .O(N__43505),
            .I(N__43490));
    LocalMux I__10059 (
            .O(N__43502),
            .I(N__43487));
    Span4Mux_h I__10058 (
            .O(N__43499),
            .I(N__43480));
    LocalMux I__10057 (
            .O(N__43496),
            .I(N__43480));
    Span4Mux_h I__10056 (
            .O(N__43493),
            .I(N__43480));
    Odrv4 I__10055 (
            .O(N__43490),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    Odrv12 I__10054 (
            .O(N__43487),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    Odrv4 I__10053 (
            .O(N__43480),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ));
    InMux I__10052 (
            .O(N__43473),
            .I(N__43455));
    InMux I__10051 (
            .O(N__43472),
            .I(N__43455));
    InMux I__10050 (
            .O(N__43471),
            .I(N__43455));
    InMux I__10049 (
            .O(N__43470),
            .I(N__43455));
    InMux I__10048 (
            .O(N__43469),
            .I(N__43455));
    InMux I__10047 (
            .O(N__43468),
            .I(N__43455));
    LocalMux I__10046 (
            .O(N__43455),
            .I(N__43439));
    InMux I__10045 (
            .O(N__43454),
            .I(N__43430));
    InMux I__10044 (
            .O(N__43453),
            .I(N__43430));
    InMux I__10043 (
            .O(N__43452),
            .I(N__43430));
    InMux I__10042 (
            .O(N__43451),
            .I(N__43430));
    InMux I__10041 (
            .O(N__43450),
            .I(N__43425));
    InMux I__10040 (
            .O(N__43449),
            .I(N__43412));
    InMux I__10039 (
            .O(N__43448),
            .I(N__43412));
    InMux I__10038 (
            .O(N__43447),
            .I(N__43412));
    InMux I__10037 (
            .O(N__43446),
            .I(N__43412));
    InMux I__10036 (
            .O(N__43445),
            .I(N__43412));
    InMux I__10035 (
            .O(N__43444),
            .I(N__43412));
    InMux I__10034 (
            .O(N__43443),
            .I(N__43407));
    InMux I__10033 (
            .O(N__43442),
            .I(N__43407));
    Span4Mux_v I__10032 (
            .O(N__43439),
            .I(N__43402));
    LocalMux I__10031 (
            .O(N__43430),
            .I(N__43402));
    InMux I__10030 (
            .O(N__43429),
            .I(N__43398));
    InMux I__10029 (
            .O(N__43428),
            .I(N__43393));
    LocalMux I__10028 (
            .O(N__43425),
            .I(N__43390));
    LocalMux I__10027 (
            .O(N__43412),
            .I(N__43387));
    LocalMux I__10026 (
            .O(N__43407),
            .I(N__43382));
    Span4Mux_h I__10025 (
            .O(N__43402),
            .I(N__43382));
    InMux I__10024 (
            .O(N__43401),
            .I(N__43379));
    LocalMux I__10023 (
            .O(N__43398),
            .I(N__43376));
    InMux I__10022 (
            .O(N__43397),
            .I(N__43373));
    InMux I__10021 (
            .O(N__43396),
            .I(N__43370));
    LocalMux I__10020 (
            .O(N__43393),
            .I(N__43363));
    Span4Mux_v I__10019 (
            .O(N__43390),
            .I(N__43363));
    Span4Mux_v I__10018 (
            .O(N__43387),
            .I(N__43363));
    Span4Mux_v I__10017 (
            .O(N__43382),
            .I(N__43358));
    LocalMux I__10016 (
            .O(N__43379),
            .I(N__43358));
    Span4Mux_h I__10015 (
            .O(N__43376),
            .I(N__43355));
    LocalMux I__10014 (
            .O(N__43373),
            .I(N__43352));
    LocalMux I__10013 (
            .O(N__43370),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10012 (
            .O(N__43363),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10011 (
            .O(N__43358),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv4 I__10010 (
            .O(N__43355),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    Odrv12 I__10009 (
            .O(N__43352),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ));
    CascadeMux I__10008 (
            .O(N__43341),
            .I(N__43327));
    CascadeMux I__10007 (
            .O(N__43340),
            .I(N__43324));
    CascadeMux I__10006 (
            .O(N__43339),
            .I(N__43321));
    CascadeMux I__10005 (
            .O(N__43338),
            .I(N__43318));
    CascadeMux I__10004 (
            .O(N__43337),
            .I(N__43312));
    CascadeMux I__10003 (
            .O(N__43336),
            .I(N__43308));
    CascadeMux I__10002 (
            .O(N__43335),
            .I(N__43305));
    CascadeMux I__10001 (
            .O(N__43334),
            .I(N__43302));
    CascadeMux I__10000 (
            .O(N__43333),
            .I(N__43299));
    CascadeMux I__9999 (
            .O(N__43332),
            .I(N__43296));
    CascadeMux I__9998 (
            .O(N__43331),
            .I(N__43293));
    InMux I__9997 (
            .O(N__43330),
            .I(N__43287));
    InMux I__9996 (
            .O(N__43327),
            .I(N__43270));
    InMux I__9995 (
            .O(N__43324),
            .I(N__43270));
    InMux I__9994 (
            .O(N__43321),
            .I(N__43270));
    InMux I__9993 (
            .O(N__43318),
            .I(N__43270));
    InMux I__9992 (
            .O(N__43317),
            .I(N__43270));
    InMux I__9991 (
            .O(N__43316),
            .I(N__43270));
    InMux I__9990 (
            .O(N__43315),
            .I(N__43265));
    InMux I__9989 (
            .O(N__43312),
            .I(N__43265));
    InMux I__9988 (
            .O(N__43311),
            .I(N__43256));
    InMux I__9987 (
            .O(N__43308),
            .I(N__43256));
    InMux I__9986 (
            .O(N__43305),
            .I(N__43256));
    InMux I__9985 (
            .O(N__43302),
            .I(N__43256));
    InMux I__9984 (
            .O(N__43299),
            .I(N__43243));
    InMux I__9983 (
            .O(N__43296),
            .I(N__43243));
    InMux I__9982 (
            .O(N__43293),
            .I(N__43243));
    InMux I__9981 (
            .O(N__43292),
            .I(N__43243));
    InMux I__9980 (
            .O(N__43291),
            .I(N__43243));
    InMux I__9979 (
            .O(N__43290),
            .I(N__43243));
    LocalMux I__9978 (
            .O(N__43287),
            .I(N__43240));
    InMux I__9977 (
            .O(N__43286),
            .I(N__43237));
    InMux I__9976 (
            .O(N__43285),
            .I(N__43234));
    CascadeMux I__9975 (
            .O(N__43284),
            .I(N__43231));
    CascadeMux I__9974 (
            .O(N__43283),
            .I(N__43228));
    LocalMux I__9973 (
            .O(N__43270),
            .I(N__43224));
    LocalMux I__9972 (
            .O(N__43265),
            .I(N__43221));
    LocalMux I__9971 (
            .O(N__43256),
            .I(N__43216));
    LocalMux I__9970 (
            .O(N__43243),
            .I(N__43216));
    Span4Mux_v I__9969 (
            .O(N__43240),
            .I(N__43211));
    LocalMux I__9968 (
            .O(N__43237),
            .I(N__43211));
    LocalMux I__9967 (
            .O(N__43234),
            .I(N__43208));
    InMux I__9966 (
            .O(N__43231),
            .I(N__43205));
    InMux I__9965 (
            .O(N__43228),
            .I(N__43200));
    InMux I__9964 (
            .O(N__43227),
            .I(N__43200));
    Span4Mux_v I__9963 (
            .O(N__43224),
            .I(N__43197));
    Span4Mux_v I__9962 (
            .O(N__43221),
            .I(N__43194));
    Span4Mux_v I__9961 (
            .O(N__43216),
            .I(N__43187));
    Span4Mux_h I__9960 (
            .O(N__43211),
            .I(N__43187));
    Span4Mux_h I__9959 (
            .O(N__43208),
            .I(N__43187));
    LocalMux I__9958 (
            .O(N__43205),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__9957 (
            .O(N__43200),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__9956 (
            .O(N__43197),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__9955 (
            .O(N__43194),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__9954 (
            .O(N__43187),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__9953 (
            .O(N__43176),
            .I(N__43173));
    LocalMux I__9952 (
            .O(N__43173),
            .I(N__43169));
    InMux I__9951 (
            .O(N__43172),
            .I(N__43166));
    Span4Mux_v I__9950 (
            .O(N__43169),
            .I(N__43160));
    LocalMux I__9949 (
            .O(N__43166),
            .I(N__43160));
    InMux I__9948 (
            .O(N__43165),
            .I(N__43157));
    Span4Mux_h I__9947 (
            .O(N__43160),
            .I(N__43152));
    LocalMux I__9946 (
            .O(N__43157),
            .I(N__43149));
    InMux I__9945 (
            .O(N__43156),
            .I(N__43146));
    InMux I__9944 (
            .O(N__43155),
            .I(N__43143));
    Span4Mux_v I__9943 (
            .O(N__43152),
            .I(N__43140));
    Span4Mux_v I__9942 (
            .O(N__43149),
            .I(N__43133));
    LocalMux I__9941 (
            .O(N__43146),
            .I(N__43133));
    LocalMux I__9940 (
            .O(N__43143),
            .I(N__43133));
    Odrv4 I__9939 (
            .O(N__43140),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9938 (
            .O(N__43133),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__9937 (
            .O(N__43128),
            .I(N__43121));
    CascadeMux I__9936 (
            .O(N__43127),
            .I(N__43118));
    CascadeMux I__9935 (
            .O(N__43126),
            .I(N__43111));
    CascadeMux I__9934 (
            .O(N__43125),
            .I(N__43105));
    CascadeMux I__9933 (
            .O(N__43124),
            .I(N__43102));
    InMux I__9932 (
            .O(N__43121),
            .I(N__43093));
    InMux I__9931 (
            .O(N__43118),
            .I(N__43093));
    InMux I__9930 (
            .O(N__43117),
            .I(N__43084));
    InMux I__9929 (
            .O(N__43116),
            .I(N__43084));
    InMux I__9928 (
            .O(N__43115),
            .I(N__43084));
    InMux I__9927 (
            .O(N__43114),
            .I(N__43084));
    InMux I__9926 (
            .O(N__43111),
            .I(N__43080));
    InMux I__9925 (
            .O(N__43110),
            .I(N__43073));
    InMux I__9924 (
            .O(N__43109),
            .I(N__43073));
    InMux I__9923 (
            .O(N__43108),
            .I(N__43073));
    InMux I__9922 (
            .O(N__43105),
            .I(N__43062));
    InMux I__9921 (
            .O(N__43102),
            .I(N__43062));
    InMux I__9920 (
            .O(N__43101),
            .I(N__43062));
    InMux I__9919 (
            .O(N__43100),
            .I(N__43055));
    InMux I__9918 (
            .O(N__43099),
            .I(N__43055));
    InMux I__9917 (
            .O(N__43098),
            .I(N__43055));
    LocalMux I__9916 (
            .O(N__43093),
            .I(N__43050));
    LocalMux I__9915 (
            .O(N__43084),
            .I(N__43050));
    InMux I__9914 (
            .O(N__43083),
            .I(N__43047));
    LocalMux I__9913 (
            .O(N__43080),
            .I(N__43043));
    LocalMux I__9912 (
            .O(N__43073),
            .I(N__43040));
    InMux I__9911 (
            .O(N__43072),
            .I(N__43035));
    InMux I__9910 (
            .O(N__43071),
            .I(N__43035));
    InMux I__9909 (
            .O(N__43070),
            .I(N__43032));
    InMux I__9908 (
            .O(N__43069),
            .I(N__43028));
    LocalMux I__9907 (
            .O(N__43062),
            .I(N__43023));
    LocalMux I__9906 (
            .O(N__43055),
            .I(N__43023));
    Span4Mux_v I__9905 (
            .O(N__43050),
            .I(N__43018));
    LocalMux I__9904 (
            .O(N__43047),
            .I(N__43018));
    InMux I__9903 (
            .O(N__43046),
            .I(N__43015));
    Span4Mux_h I__9902 (
            .O(N__43043),
            .I(N__43006));
    Span4Mux_h I__9901 (
            .O(N__43040),
            .I(N__43006));
    LocalMux I__9900 (
            .O(N__43035),
            .I(N__43006));
    LocalMux I__9899 (
            .O(N__43032),
            .I(N__43006));
    CascadeMux I__9898 (
            .O(N__43031),
            .I(N__43003));
    LocalMux I__9897 (
            .O(N__43028),
            .I(N__43000));
    Span4Mux_h I__9896 (
            .O(N__43023),
            .I(N__42997));
    Span4Mux_v I__9895 (
            .O(N__43018),
            .I(N__42993));
    LocalMux I__9894 (
            .O(N__43015),
            .I(N__42988));
    Span4Mux_v I__9893 (
            .O(N__43006),
            .I(N__42988));
    InMux I__9892 (
            .O(N__43003),
            .I(N__42985));
    Span4Mux_v I__9891 (
            .O(N__43000),
            .I(N__42982));
    Span4Mux_v I__9890 (
            .O(N__42997),
            .I(N__42979));
    InMux I__9889 (
            .O(N__42996),
            .I(N__42976));
    Span4Mux_h I__9888 (
            .O(N__42993),
            .I(N__42971));
    Span4Mux_v I__9887 (
            .O(N__42988),
            .I(N__42971));
    LocalMux I__9886 (
            .O(N__42985),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9885 (
            .O(N__42982),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9884 (
            .O(N__42979),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    LocalMux I__9883 (
            .O(N__42976),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    Odrv4 I__9882 (
            .O(N__42971),
            .I(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ));
    CascadeMux I__9881 (
            .O(N__42960),
            .I(N__42944));
    CascadeMux I__9880 (
            .O(N__42959),
            .I(N__42940));
    CascadeMux I__9879 (
            .O(N__42958),
            .I(N__42931));
    CascadeMux I__9878 (
            .O(N__42957),
            .I(N__42928));
    CascadeMux I__9877 (
            .O(N__42956),
            .I(N__42925));
    CascadeMux I__9876 (
            .O(N__42955),
            .I(N__42922));
    CascadeMux I__9875 (
            .O(N__42954),
            .I(N__42919));
    InMux I__9874 (
            .O(N__42953),
            .I(N__42905));
    InMux I__9873 (
            .O(N__42952),
            .I(N__42905));
    InMux I__9872 (
            .O(N__42951),
            .I(N__42905));
    InMux I__9871 (
            .O(N__42950),
            .I(N__42905));
    InMux I__9870 (
            .O(N__42949),
            .I(N__42905));
    InMux I__9869 (
            .O(N__42948),
            .I(N__42905));
    InMux I__9868 (
            .O(N__42947),
            .I(N__42902));
    InMux I__9867 (
            .O(N__42944),
            .I(N__42899));
    InMux I__9866 (
            .O(N__42943),
            .I(N__42896));
    InMux I__9865 (
            .O(N__42940),
            .I(N__42889));
    InMux I__9864 (
            .O(N__42939),
            .I(N__42889));
    InMux I__9863 (
            .O(N__42938),
            .I(N__42889));
    InMux I__9862 (
            .O(N__42937),
            .I(N__42872));
    InMux I__9861 (
            .O(N__42936),
            .I(N__42872));
    InMux I__9860 (
            .O(N__42935),
            .I(N__42872));
    InMux I__9859 (
            .O(N__42934),
            .I(N__42872));
    InMux I__9858 (
            .O(N__42931),
            .I(N__42872));
    InMux I__9857 (
            .O(N__42928),
            .I(N__42872));
    InMux I__9856 (
            .O(N__42925),
            .I(N__42872));
    InMux I__9855 (
            .O(N__42922),
            .I(N__42872));
    InMux I__9854 (
            .O(N__42919),
            .I(N__42867));
    InMux I__9853 (
            .O(N__42918),
            .I(N__42867));
    LocalMux I__9852 (
            .O(N__42905),
            .I(N__42864));
    LocalMux I__9851 (
            .O(N__42902),
            .I(N__42859));
    LocalMux I__9850 (
            .O(N__42899),
            .I(N__42859));
    LocalMux I__9849 (
            .O(N__42896),
            .I(N__42856));
    LocalMux I__9848 (
            .O(N__42889),
            .I(N__42853));
    LocalMux I__9847 (
            .O(N__42872),
            .I(N__42850));
    LocalMux I__9846 (
            .O(N__42867),
            .I(N__42839));
    Span4Mux_h I__9845 (
            .O(N__42864),
            .I(N__42839));
    Span4Mux_v I__9844 (
            .O(N__42859),
            .I(N__42839));
    Span4Mux_v I__9843 (
            .O(N__42856),
            .I(N__42839));
    Span4Mux_h I__9842 (
            .O(N__42853),
            .I(N__42834));
    Span4Mux_h I__9841 (
            .O(N__42850),
            .I(N__42834));
    InMux I__9840 (
            .O(N__42849),
            .I(N__42831));
    InMux I__9839 (
            .O(N__42848),
            .I(N__42828));
    Odrv4 I__9838 (
            .O(N__42839),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__9837 (
            .O(N__42834),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__9836 (
            .O(N__42831),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__9835 (
            .O(N__42828),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__9834 (
            .O(N__42819),
            .I(N__42816));
    InMux I__9833 (
            .O(N__42816),
            .I(N__42809));
    InMux I__9832 (
            .O(N__42815),
            .I(N__42798));
    InMux I__9831 (
            .O(N__42814),
            .I(N__42798));
    InMux I__9830 (
            .O(N__42813),
            .I(N__42798));
    InMux I__9829 (
            .O(N__42812),
            .I(N__42794));
    LocalMux I__9828 (
            .O(N__42809),
            .I(N__42782));
    CascadeMux I__9827 (
            .O(N__42808),
            .I(N__42777));
    CascadeMux I__9826 (
            .O(N__42807),
            .I(N__42772));
    CascadeMux I__9825 (
            .O(N__42806),
            .I(N__42769));
    CascadeMux I__9824 (
            .O(N__42805),
            .I(N__42766));
    LocalMux I__9823 (
            .O(N__42798),
            .I(N__42763));
    InMux I__9822 (
            .O(N__42797),
            .I(N__42760));
    LocalMux I__9821 (
            .O(N__42794),
            .I(N__42757));
    InMux I__9820 (
            .O(N__42793),
            .I(N__42754));
    InMux I__9819 (
            .O(N__42792),
            .I(N__42736));
    InMux I__9818 (
            .O(N__42791),
            .I(N__42736));
    InMux I__9817 (
            .O(N__42790),
            .I(N__42736));
    InMux I__9816 (
            .O(N__42789),
            .I(N__42736));
    InMux I__9815 (
            .O(N__42788),
            .I(N__42736));
    InMux I__9814 (
            .O(N__42787),
            .I(N__42736));
    InMux I__9813 (
            .O(N__42786),
            .I(N__42736));
    InMux I__9812 (
            .O(N__42785),
            .I(N__42736));
    Span4Mux_v I__9811 (
            .O(N__42782),
            .I(N__42733));
    InMux I__9810 (
            .O(N__42781),
            .I(N__42730));
    InMux I__9809 (
            .O(N__42780),
            .I(N__42725));
    InMux I__9808 (
            .O(N__42777),
            .I(N__42725));
    InMux I__9807 (
            .O(N__42776),
            .I(N__42714));
    InMux I__9806 (
            .O(N__42775),
            .I(N__42714));
    InMux I__9805 (
            .O(N__42772),
            .I(N__42714));
    InMux I__9804 (
            .O(N__42769),
            .I(N__42714));
    InMux I__9803 (
            .O(N__42766),
            .I(N__42714));
    Span4Mux_v I__9802 (
            .O(N__42763),
            .I(N__42711));
    LocalMux I__9801 (
            .O(N__42760),
            .I(N__42704));
    Span4Mux_v I__9800 (
            .O(N__42757),
            .I(N__42704));
    LocalMux I__9799 (
            .O(N__42754),
            .I(N__42704));
    InMux I__9798 (
            .O(N__42753),
            .I(N__42701));
    LocalMux I__9797 (
            .O(N__42736),
            .I(N__42694));
    Span4Mux_h I__9796 (
            .O(N__42733),
            .I(N__42694));
    LocalMux I__9795 (
            .O(N__42730),
            .I(N__42694));
    LocalMux I__9794 (
            .O(N__42725),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__9793 (
            .O(N__42714),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__9792 (
            .O(N__42711),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__9791 (
            .O(N__42704),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__9790 (
            .O(N__42701),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__9789 (
            .O(N__42694),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ));
    InMux I__9788 (
            .O(N__42681),
            .I(N__42677));
    InMux I__9787 (
            .O(N__42680),
            .I(N__42674));
    LocalMux I__9786 (
            .O(N__42677),
            .I(N__42669));
    LocalMux I__9785 (
            .O(N__42674),
            .I(N__42666));
    InMux I__9784 (
            .O(N__42673),
            .I(N__42663));
    InMux I__9783 (
            .O(N__42672),
            .I(N__42660));
    Span4Mux_v I__9782 (
            .O(N__42669),
            .I(N__42655));
    Span12Mux_v I__9781 (
            .O(N__42666),
            .I(N__42652));
    LocalMux I__9780 (
            .O(N__42663),
            .I(N__42649));
    LocalMux I__9779 (
            .O(N__42660),
            .I(N__42646));
    InMux I__9778 (
            .O(N__42659),
            .I(N__42641));
    InMux I__9777 (
            .O(N__42658),
            .I(N__42641));
    Odrv4 I__9776 (
            .O(N__42655),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv12 I__9775 (
            .O(N__42652),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9774 (
            .O(N__42649),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__9773 (
            .O(N__42646),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    LocalMux I__9772 (
            .O(N__42641),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    InMux I__9771 (
            .O(N__42630),
            .I(N__42614));
    InMux I__9770 (
            .O(N__42629),
            .I(N__42611));
    InMux I__9769 (
            .O(N__42628),
            .I(N__42600));
    InMux I__9768 (
            .O(N__42627),
            .I(N__42585));
    InMux I__9767 (
            .O(N__42626),
            .I(N__42585));
    InMux I__9766 (
            .O(N__42625),
            .I(N__42585));
    InMux I__9765 (
            .O(N__42624),
            .I(N__42585));
    InMux I__9764 (
            .O(N__42623),
            .I(N__42585));
    InMux I__9763 (
            .O(N__42622),
            .I(N__42585));
    InMux I__9762 (
            .O(N__42621),
            .I(N__42585));
    InMux I__9761 (
            .O(N__42620),
            .I(N__42582));
    InMux I__9760 (
            .O(N__42619),
            .I(N__42574));
    InMux I__9759 (
            .O(N__42618),
            .I(N__42574));
    InMux I__9758 (
            .O(N__42617),
            .I(N__42574));
    LocalMux I__9757 (
            .O(N__42614),
            .I(N__42569));
    LocalMux I__9756 (
            .O(N__42611),
            .I(N__42569));
    InMux I__9755 (
            .O(N__42610),
            .I(N__42552));
    InMux I__9754 (
            .O(N__42609),
            .I(N__42552));
    InMux I__9753 (
            .O(N__42608),
            .I(N__42552));
    InMux I__9752 (
            .O(N__42607),
            .I(N__42552));
    InMux I__9751 (
            .O(N__42606),
            .I(N__42552));
    InMux I__9750 (
            .O(N__42605),
            .I(N__42552));
    InMux I__9749 (
            .O(N__42604),
            .I(N__42552));
    InMux I__9748 (
            .O(N__42603),
            .I(N__42552));
    LocalMux I__9747 (
            .O(N__42600),
            .I(N__42549));
    LocalMux I__9746 (
            .O(N__42585),
            .I(N__42544));
    LocalMux I__9745 (
            .O(N__42582),
            .I(N__42544));
    InMux I__9744 (
            .O(N__42581),
            .I(N__42541));
    LocalMux I__9743 (
            .O(N__42574),
            .I(N__42535));
    Span4Mux_h I__9742 (
            .O(N__42569),
            .I(N__42535));
    LocalMux I__9741 (
            .O(N__42552),
            .I(N__42526));
    Span4Mux_h I__9740 (
            .O(N__42549),
            .I(N__42526));
    Span4Mux_v I__9739 (
            .O(N__42544),
            .I(N__42526));
    LocalMux I__9738 (
            .O(N__42541),
            .I(N__42526));
    InMux I__9737 (
            .O(N__42540),
            .I(N__42523));
    Span4Mux_v I__9736 (
            .O(N__42535),
            .I(N__42520));
    Span4Mux_v I__9735 (
            .O(N__42526),
            .I(N__42517));
    LocalMux I__9734 (
            .O(N__42523),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__9733 (
            .O(N__42520),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__9732 (
            .O(N__42517),
            .I(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ));
    CEMux I__9731 (
            .O(N__42510),
            .I(N__42503));
    CEMux I__9730 (
            .O(N__42509),
            .I(N__42499));
    CEMux I__9729 (
            .O(N__42508),
            .I(N__42496));
    CEMux I__9728 (
            .O(N__42507),
            .I(N__42493));
    IoInMux I__9727 (
            .O(N__42506),
            .I(N__42490));
    LocalMux I__9726 (
            .O(N__42503),
            .I(N__42487));
    CEMux I__9725 (
            .O(N__42502),
            .I(N__42484));
    LocalMux I__9724 (
            .O(N__42499),
            .I(N__42481));
    LocalMux I__9723 (
            .O(N__42496),
            .I(N__42478));
    LocalMux I__9722 (
            .O(N__42493),
            .I(N__42475));
    LocalMux I__9721 (
            .O(N__42490),
            .I(N__42472));
    Span4Mux_v I__9720 (
            .O(N__42487),
            .I(N__42469));
    LocalMux I__9719 (
            .O(N__42484),
            .I(N__42466));
    Span12Mux_h I__9718 (
            .O(N__42481),
            .I(N__42463));
    Span12Mux_s10_v I__9717 (
            .O(N__42478),
            .I(N__42458));
    Sp12to4 I__9716 (
            .O(N__42475),
            .I(N__42458));
    Span4Mux_s3_v I__9715 (
            .O(N__42472),
            .I(N__42455));
    Span4Mux_v I__9714 (
            .O(N__42469),
            .I(N__42452));
    Span4Mux_v I__9713 (
            .O(N__42466),
            .I(N__42449));
    Span12Mux_v I__9712 (
            .O(N__42463),
            .I(N__42446));
    Span12Mux_v I__9711 (
            .O(N__42458),
            .I(N__42443));
    Span4Mux_v I__9710 (
            .O(N__42455),
            .I(N__42440));
    Span4Mux_v I__9709 (
            .O(N__42452),
            .I(N__42437));
    Span4Mux_v I__9708 (
            .O(N__42449),
            .I(N__42434));
    Odrv12 I__9707 (
            .O(N__42446),
            .I(red_c_i));
    Odrv12 I__9706 (
            .O(N__42443),
            .I(red_c_i));
    Odrv4 I__9705 (
            .O(N__42440),
            .I(red_c_i));
    Odrv4 I__9704 (
            .O(N__42437),
            .I(red_c_i));
    Odrv4 I__9703 (
            .O(N__42434),
            .I(red_c_i));
    InMux I__9702 (
            .O(N__42423),
            .I(N__42419));
    InMux I__9701 (
            .O(N__42422),
            .I(N__42416));
    LocalMux I__9700 (
            .O(N__42419),
            .I(N__42411));
    LocalMux I__9699 (
            .O(N__42416),
            .I(N__42411));
    Span4Mux_v I__9698 (
            .O(N__42411),
            .I(N__42408));
    Odrv4 I__9697 (
            .O(N__42408),
            .I(\delay_measurement_inst.elapsed_time_hc_1 ));
    CascadeMux I__9696 (
            .O(N__42405),
            .I(N__42402));
    InMux I__9695 (
            .O(N__42402),
            .I(N__42397));
    InMux I__9694 (
            .O(N__42401),
            .I(N__42394));
    CascadeMux I__9693 (
            .O(N__42400),
            .I(N__42391));
    LocalMux I__9692 (
            .O(N__42397),
            .I(N__42388));
    LocalMux I__9691 (
            .O(N__42394),
            .I(N__42385));
    InMux I__9690 (
            .O(N__42391),
            .I(N__42382));
    Span4Mux_h I__9689 (
            .O(N__42388),
            .I(N__42379));
    Odrv4 I__9688 (
            .O(N__42385),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    LocalMux I__9687 (
            .O(N__42382),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    Odrv4 I__9686 (
            .O(N__42379),
            .I(\delay_measurement_inst.elapsed_time_hc_3 ));
    InMux I__9685 (
            .O(N__42372),
            .I(N__42368));
    InMux I__9684 (
            .O(N__42371),
            .I(N__42365));
    LocalMux I__9683 (
            .O(N__42368),
            .I(N__42362));
    LocalMux I__9682 (
            .O(N__42365),
            .I(N__42359));
    Span4Mux_v I__9681 (
            .O(N__42362),
            .I(N__42353));
    Span4Mux_h I__9680 (
            .O(N__42359),
            .I(N__42353));
    InMux I__9679 (
            .O(N__42358),
            .I(N__42350));
    Odrv4 I__9678 (
            .O(N__42353),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    LocalMux I__9677 (
            .O(N__42350),
            .I(\delay_measurement_inst.elapsed_time_hc_5 ));
    InMux I__9676 (
            .O(N__42345),
            .I(N__42342));
    LocalMux I__9675 (
            .O(N__42342),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_3 ));
    InMux I__9674 (
            .O(N__42339),
            .I(N__42336));
    LocalMux I__9673 (
            .O(N__42336),
            .I(N__42332));
    InMux I__9672 (
            .O(N__42335),
            .I(N__42329));
    Span4Mux_v I__9671 (
            .O(N__42332),
            .I(N__42326));
    LocalMux I__9670 (
            .O(N__42329),
            .I(N__42323));
    Odrv4 I__9669 (
            .O(N__42326),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    Odrv4 I__9668 (
            .O(N__42323),
            .I(\delay_measurement_inst.delay_hc_reg3lto6 ));
    InMux I__9667 (
            .O(N__42318),
            .I(N__42314));
    InMux I__9666 (
            .O(N__42317),
            .I(N__42311));
    LocalMux I__9665 (
            .O(N__42314),
            .I(\delay_measurement_inst.N_332 ));
    LocalMux I__9664 (
            .O(N__42311),
            .I(\delay_measurement_inst.N_332 ));
    InMux I__9663 (
            .O(N__42306),
            .I(N__42302));
    InMux I__9662 (
            .O(N__42305),
            .I(N__42299));
    LocalMux I__9661 (
            .O(N__42302),
            .I(\delay_measurement_inst.N_318 ));
    LocalMux I__9660 (
            .O(N__42299),
            .I(\delay_measurement_inst.N_318 ));
    InMux I__9659 (
            .O(N__42294),
            .I(N__42291));
    LocalMux I__9658 (
            .O(N__42291),
            .I(N__42288));
    Odrv12 I__9657 (
            .O(N__42288),
            .I(\delay_measurement_inst.N_295 ));
    InMux I__9656 (
            .O(N__42285),
            .I(N__42282));
    LocalMux I__9655 (
            .O(N__42282),
            .I(N__42279));
    Span4Mux_h I__9654 (
            .O(N__42279),
            .I(N__42273));
    InMux I__9653 (
            .O(N__42278),
            .I(N__42266));
    InMux I__9652 (
            .O(N__42277),
            .I(N__42266));
    InMux I__9651 (
            .O(N__42276),
            .I(N__42266));
    Odrv4 I__9650 (
            .O(N__42273),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    LocalMux I__9649 (
            .O(N__42266),
            .I(\delay_measurement_inst.delay_hc_reg3lto15 ));
    InMux I__9648 (
            .O(N__42261),
            .I(N__42253));
    InMux I__9647 (
            .O(N__42260),
            .I(N__42250));
    InMux I__9646 (
            .O(N__42259),
            .I(N__42247));
    InMux I__9645 (
            .O(N__42258),
            .I(N__42242));
    InMux I__9644 (
            .O(N__42257),
            .I(N__42242));
    CascadeMux I__9643 (
            .O(N__42256),
            .I(N__42239));
    LocalMux I__9642 (
            .O(N__42253),
            .I(N__42232));
    LocalMux I__9641 (
            .O(N__42250),
            .I(N__42232));
    LocalMux I__9640 (
            .O(N__42247),
            .I(N__42232));
    LocalMux I__9639 (
            .O(N__42242),
            .I(N__42229));
    InMux I__9638 (
            .O(N__42239),
            .I(N__42226));
    Sp12to4 I__9637 (
            .O(N__42232),
            .I(N__42223));
    Span4Mux_h I__9636 (
            .O(N__42229),
            .I(N__42220));
    LocalMux I__9635 (
            .O(N__42226),
            .I(measured_delay_hc_15));
    Odrv12 I__9634 (
            .O(N__42223),
            .I(measured_delay_hc_15));
    Odrv4 I__9633 (
            .O(N__42220),
            .I(measured_delay_hc_15));
    CascadeMux I__9632 (
            .O(N__42213),
            .I(N__42210));
    InMux I__9631 (
            .O(N__42210),
            .I(N__42207));
    LocalMux I__9630 (
            .O(N__42207),
            .I(N__42204));
    Span4Mux_h I__9629 (
            .O(N__42204),
            .I(N__42201));
    Odrv4 I__9628 (
            .O(N__42201),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ));
    InMux I__9627 (
            .O(N__42198),
            .I(N__42194));
    InMux I__9626 (
            .O(N__42197),
            .I(N__42191));
    LocalMux I__9625 (
            .O(N__42194),
            .I(N__42188));
    LocalMux I__9624 (
            .O(N__42191),
            .I(N__42185));
    Span4Mux_v I__9623 (
            .O(N__42188),
            .I(N__42182));
    Span4Mux_v I__9622 (
            .O(N__42185),
            .I(N__42179));
    Span4Mux_h I__9621 (
            .O(N__42182),
            .I(N__42176));
    Span4Mux_h I__9620 (
            .O(N__42179),
            .I(N__42173));
    Odrv4 I__9619 (
            .O(N__42176),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__9618 (
            .O(N__42173),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__9617 (
            .O(N__42168),
            .I(N__42165));
    LocalMux I__9616 (
            .O(N__42165),
            .I(N__42162));
    Span4Mux_h I__9615 (
            .O(N__42162),
            .I(N__42159));
    Odrv4 I__9614 (
            .O(N__42159),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ));
    InMux I__9613 (
            .O(N__42156),
            .I(N__42152));
    InMux I__9612 (
            .O(N__42155),
            .I(N__42149));
    LocalMux I__9611 (
            .O(N__42152),
            .I(N__42146));
    LocalMux I__9610 (
            .O(N__42149),
            .I(N__42143));
    Span4Mux_v I__9609 (
            .O(N__42146),
            .I(N__42140));
    Span12Mux_s8_v I__9608 (
            .O(N__42143),
            .I(N__42137));
    Odrv4 I__9607 (
            .O(N__42140),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__9606 (
            .O(N__42137),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__9605 (
            .O(N__42132),
            .I(N__42129));
    InMux I__9604 (
            .O(N__42129),
            .I(N__42126));
    LocalMux I__9603 (
            .O(N__42126),
            .I(N__42123));
    Odrv12 I__9602 (
            .O(N__42123),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ));
    InMux I__9601 (
            .O(N__42120),
            .I(N__42116));
    InMux I__9600 (
            .O(N__42119),
            .I(N__42113));
    LocalMux I__9599 (
            .O(N__42116),
            .I(N__42108));
    LocalMux I__9598 (
            .O(N__42113),
            .I(N__42108));
    Odrv12 I__9597 (
            .O(N__42108),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__9596 (
            .O(N__42105),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__9595 (
            .O(N__42102),
            .I(N__42098));
    InMux I__9594 (
            .O(N__42101),
            .I(N__42095));
    LocalMux I__9593 (
            .O(N__42098),
            .I(measured_delay_hc_27));
    LocalMux I__9592 (
            .O(N__42095),
            .I(measured_delay_hc_27));
    InMux I__9591 (
            .O(N__42090),
            .I(N__42086));
    InMux I__9590 (
            .O(N__42089),
            .I(N__42083));
    LocalMux I__9589 (
            .O(N__42086),
            .I(measured_delay_hc_28));
    LocalMux I__9588 (
            .O(N__42083),
            .I(measured_delay_hc_28));
    InMux I__9587 (
            .O(N__42078),
            .I(N__42073));
    InMux I__9586 (
            .O(N__42077),
            .I(N__42070));
    InMux I__9585 (
            .O(N__42076),
            .I(N__42067));
    LocalMux I__9584 (
            .O(N__42073),
            .I(N__42063));
    LocalMux I__9583 (
            .O(N__42070),
            .I(N__42058));
    LocalMux I__9582 (
            .O(N__42067),
            .I(N__42058));
    InMux I__9581 (
            .O(N__42066),
            .I(N__42055));
    Span4Mux_h I__9580 (
            .O(N__42063),
            .I(N__42050));
    Span4Mux_v I__9579 (
            .O(N__42058),
            .I(N__42050));
    LocalMux I__9578 (
            .O(N__42055),
            .I(measured_delay_hc_0));
    Odrv4 I__9577 (
            .O(N__42050),
            .I(measured_delay_hc_0));
    InMux I__9576 (
            .O(N__42045),
            .I(N__42041));
    CascadeMux I__9575 (
            .O(N__42044),
            .I(N__42037));
    LocalMux I__9574 (
            .O(N__42041),
            .I(N__42034));
    InMux I__9573 (
            .O(N__42040),
            .I(N__42031));
    InMux I__9572 (
            .O(N__42037),
            .I(N__42028));
    Span4Mux_v I__9571 (
            .O(N__42034),
            .I(N__42025));
    LocalMux I__9570 (
            .O(N__42031),
            .I(N__42022));
    LocalMux I__9569 (
            .O(N__42028),
            .I(N__42019));
    Span4Mux_h I__9568 (
            .O(N__42025),
            .I(N__42014));
    Span4Mux_v I__9567 (
            .O(N__42022),
            .I(N__42014));
    Span4Mux_h I__9566 (
            .O(N__42019),
            .I(N__42011));
    Odrv4 I__9565 (
            .O(N__42014),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    Odrv4 I__9564 (
            .O(N__42011),
            .I(\delay_measurement_inst.elapsed_time_hc_19 ));
    CascadeMux I__9563 (
            .O(N__42006),
            .I(N__42002));
    CascadeMux I__9562 (
            .O(N__42005),
            .I(N__41999));
    InMux I__9561 (
            .O(N__42002),
            .I(N__41994));
    InMux I__9560 (
            .O(N__41999),
            .I(N__41991));
    CascadeMux I__9559 (
            .O(N__41998),
            .I(N__41987));
    InMux I__9558 (
            .O(N__41997),
            .I(N__41984));
    LocalMux I__9557 (
            .O(N__41994),
            .I(N__41981));
    LocalMux I__9556 (
            .O(N__41991),
            .I(N__41978));
    InMux I__9555 (
            .O(N__41990),
            .I(N__41975));
    InMux I__9554 (
            .O(N__41987),
            .I(N__41972));
    LocalMux I__9553 (
            .O(N__41984),
            .I(measured_delay_hc_19));
    Odrv12 I__9552 (
            .O(N__41981),
            .I(measured_delay_hc_19));
    Odrv4 I__9551 (
            .O(N__41978),
            .I(measured_delay_hc_19));
    LocalMux I__9550 (
            .O(N__41975),
            .I(measured_delay_hc_19));
    LocalMux I__9549 (
            .O(N__41972),
            .I(measured_delay_hc_19));
    InMux I__9548 (
            .O(N__41961),
            .I(N__41958));
    LocalMux I__9547 (
            .O(N__41958),
            .I(N__41955));
    Span4Mux_h I__9546 (
            .O(N__41955),
            .I(N__41950));
    InMux I__9545 (
            .O(N__41954),
            .I(N__41945));
    InMux I__9544 (
            .O(N__41953),
            .I(N__41945));
    Odrv4 I__9543 (
            .O(N__41950),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    LocalMux I__9542 (
            .O(N__41945),
            .I(\delay_measurement_inst.elapsed_time_hc_16 ));
    InMux I__9541 (
            .O(N__41940),
            .I(N__41937));
    LocalMux I__9540 (
            .O(N__41937),
            .I(N__41931));
    InMux I__9539 (
            .O(N__41936),
            .I(N__41928));
    InMux I__9538 (
            .O(N__41935),
            .I(N__41925));
    InMux I__9537 (
            .O(N__41934),
            .I(N__41922));
    Span4Mux_h I__9536 (
            .O(N__41931),
            .I(N__41918));
    LocalMux I__9535 (
            .O(N__41928),
            .I(N__41911));
    LocalMux I__9534 (
            .O(N__41925),
            .I(N__41911));
    LocalMux I__9533 (
            .O(N__41922),
            .I(N__41911));
    InMux I__9532 (
            .O(N__41921),
            .I(N__41908));
    Span4Mux_v I__9531 (
            .O(N__41918),
            .I(N__41905));
    Span4Mux_v I__9530 (
            .O(N__41911),
            .I(N__41902));
    LocalMux I__9529 (
            .O(N__41908),
            .I(measured_delay_hc_1));
    Odrv4 I__9528 (
            .O(N__41905),
            .I(measured_delay_hc_1));
    Odrv4 I__9527 (
            .O(N__41902),
            .I(measured_delay_hc_1));
    CascadeMux I__9526 (
            .O(N__41895),
            .I(N__41892));
    InMux I__9525 (
            .O(N__41892),
            .I(N__41889));
    LocalMux I__9524 (
            .O(N__41889),
            .I(N__41886));
    Span4Mux_h I__9523 (
            .O(N__41886),
            .I(N__41881));
    InMux I__9522 (
            .O(N__41885),
            .I(N__41878));
    InMux I__9521 (
            .O(N__41884),
            .I(N__41875));
    Odrv4 I__9520 (
            .O(N__41881),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__9519 (
            .O(N__41878),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    LocalMux I__9518 (
            .O(N__41875),
            .I(\delay_measurement_inst.elapsed_time_hc_18 ));
    InMux I__9517 (
            .O(N__41868),
            .I(N__41863));
    InMux I__9516 (
            .O(N__41867),
            .I(N__41860));
    InMux I__9515 (
            .O(N__41866),
            .I(N__41855));
    LocalMux I__9514 (
            .O(N__41863),
            .I(N__41850));
    LocalMux I__9513 (
            .O(N__41860),
            .I(N__41850));
    InMux I__9512 (
            .O(N__41859),
            .I(N__41847));
    InMux I__9511 (
            .O(N__41858),
            .I(N__41844));
    LocalMux I__9510 (
            .O(N__41855),
            .I(N__41841));
    Span4Mux_v I__9509 (
            .O(N__41850),
            .I(N__41836));
    LocalMux I__9508 (
            .O(N__41847),
            .I(N__41836));
    LocalMux I__9507 (
            .O(N__41844),
            .I(measured_delay_hc_18));
    Odrv4 I__9506 (
            .O(N__41841),
            .I(measured_delay_hc_18));
    Odrv4 I__9505 (
            .O(N__41836),
            .I(measured_delay_hc_18));
    InMux I__9504 (
            .O(N__41829),
            .I(N__41824));
    InMux I__9503 (
            .O(N__41828),
            .I(N__41821));
    CascadeMux I__9502 (
            .O(N__41827),
            .I(N__41818));
    LocalMux I__9501 (
            .O(N__41824),
            .I(N__41811));
    LocalMux I__9500 (
            .O(N__41821),
            .I(N__41811));
    InMux I__9499 (
            .O(N__41818),
            .I(N__41808));
    CascadeMux I__9498 (
            .O(N__41817),
            .I(N__41805));
    InMux I__9497 (
            .O(N__41816),
            .I(N__41802));
    Span4Mux_v I__9496 (
            .O(N__41811),
            .I(N__41797));
    LocalMux I__9495 (
            .O(N__41808),
            .I(N__41797));
    InMux I__9494 (
            .O(N__41805),
            .I(N__41794));
    LocalMux I__9493 (
            .O(N__41802),
            .I(N__41791));
    Span4Mux_h I__9492 (
            .O(N__41797),
            .I(N__41788));
    LocalMux I__9491 (
            .O(N__41794),
            .I(measured_delay_hc_13));
    Odrv4 I__9490 (
            .O(N__41791),
            .I(measured_delay_hc_13));
    Odrv4 I__9489 (
            .O(N__41788),
            .I(measured_delay_hc_13));
    CascadeMux I__9488 (
            .O(N__41781),
            .I(N__41775));
    CascadeMux I__9487 (
            .O(N__41780),
            .I(N__41772));
    CascadeMux I__9486 (
            .O(N__41779),
            .I(N__41765));
    InMux I__9485 (
            .O(N__41778),
            .I(N__41754));
    InMux I__9484 (
            .O(N__41775),
            .I(N__41754));
    InMux I__9483 (
            .O(N__41772),
            .I(N__41754));
    InMux I__9482 (
            .O(N__41771),
            .I(N__41754));
    CascadeMux I__9481 (
            .O(N__41770),
            .I(N__41743));
    CascadeMux I__9480 (
            .O(N__41769),
            .I(N__41740));
    CascadeMux I__9479 (
            .O(N__41768),
            .I(N__41737));
    InMux I__9478 (
            .O(N__41765),
            .I(N__41726));
    InMux I__9477 (
            .O(N__41764),
            .I(N__41726));
    InMux I__9476 (
            .O(N__41763),
            .I(N__41726));
    LocalMux I__9475 (
            .O(N__41754),
            .I(N__41723));
    InMux I__9474 (
            .O(N__41753),
            .I(N__41708));
    InMux I__9473 (
            .O(N__41752),
            .I(N__41708));
    InMux I__9472 (
            .O(N__41751),
            .I(N__41708));
    InMux I__9471 (
            .O(N__41750),
            .I(N__41708));
    InMux I__9470 (
            .O(N__41749),
            .I(N__41708));
    InMux I__9469 (
            .O(N__41748),
            .I(N__41708));
    InMux I__9468 (
            .O(N__41747),
            .I(N__41708));
    InMux I__9467 (
            .O(N__41746),
            .I(N__41699));
    InMux I__9466 (
            .O(N__41743),
            .I(N__41699));
    InMux I__9465 (
            .O(N__41740),
            .I(N__41699));
    InMux I__9464 (
            .O(N__41737),
            .I(N__41699));
    InMux I__9463 (
            .O(N__41736),
            .I(N__41690));
    InMux I__9462 (
            .O(N__41735),
            .I(N__41690));
    InMux I__9461 (
            .O(N__41734),
            .I(N__41690));
    InMux I__9460 (
            .O(N__41733),
            .I(N__41690));
    LocalMux I__9459 (
            .O(N__41726),
            .I(N__41687));
    Span4Mux_h I__9458 (
            .O(N__41723),
            .I(N__41684));
    LocalMux I__9457 (
            .O(N__41708),
            .I(N__41681));
    LocalMux I__9456 (
            .O(N__41699),
            .I(\phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ));
    LocalMux I__9455 (
            .O(N__41690),
            .I(\phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ));
    Odrv4 I__9454 (
            .O(N__41687),
            .I(\phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ));
    Odrv4 I__9453 (
            .O(N__41684),
            .I(\phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ));
    Odrv12 I__9452 (
            .O(N__41681),
            .I(\phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ));
    InMux I__9451 (
            .O(N__41670),
            .I(N__41665));
    InMux I__9450 (
            .O(N__41669),
            .I(N__41660));
    InMux I__9449 (
            .O(N__41668),
            .I(N__41660));
    LocalMux I__9448 (
            .O(N__41665),
            .I(\phase_controller_inst1.stoper_hc.N_459 ));
    LocalMux I__9447 (
            .O(N__41660),
            .I(\phase_controller_inst1.stoper_hc.N_459 ));
    CascadeMux I__9446 (
            .O(N__41655),
            .I(N__41652));
    InMux I__9445 (
            .O(N__41652),
            .I(N__41649));
    LocalMux I__9444 (
            .O(N__41649),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3 ));
    InMux I__9443 (
            .O(N__41646),
            .I(N__41641));
    InMux I__9442 (
            .O(N__41645),
            .I(N__41638));
    InMux I__9441 (
            .O(N__41644),
            .I(N__41634));
    LocalMux I__9440 (
            .O(N__41641),
            .I(N__41629));
    LocalMux I__9439 (
            .O(N__41638),
            .I(N__41629));
    InMux I__9438 (
            .O(N__41637),
            .I(N__41626));
    LocalMux I__9437 (
            .O(N__41634),
            .I(N__41623));
    Span4Mux_v I__9436 (
            .O(N__41629),
            .I(N__41617));
    LocalMux I__9435 (
            .O(N__41626),
            .I(N__41617));
    Span4Mux_v I__9434 (
            .O(N__41623),
            .I(N__41614));
    InMux I__9433 (
            .O(N__41622),
            .I(N__41611));
    Span4Mux_h I__9432 (
            .O(N__41617),
            .I(N__41608));
    Span4Mux_h I__9431 (
            .O(N__41614),
            .I(N__41605));
    LocalMux I__9430 (
            .O(N__41611),
            .I(measured_delay_hc_3));
    Odrv4 I__9429 (
            .O(N__41608),
            .I(measured_delay_hc_3));
    Odrv4 I__9428 (
            .O(N__41605),
            .I(measured_delay_hc_3));
    CascadeMux I__9427 (
            .O(N__41598),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3_cascade_ ));
    CascadeMux I__9426 (
            .O(N__41595),
            .I(N__41589));
    CascadeMux I__9425 (
            .O(N__41594),
            .I(N__41586));
    CascadeMux I__9424 (
            .O(N__41593),
            .I(N__41583));
    CascadeMux I__9423 (
            .O(N__41592),
            .I(N__41579));
    InMux I__9422 (
            .O(N__41589),
            .I(N__41576));
    InMux I__9421 (
            .O(N__41586),
            .I(N__41573));
    InMux I__9420 (
            .O(N__41583),
            .I(N__41570));
    InMux I__9419 (
            .O(N__41582),
            .I(N__41567));
    InMux I__9418 (
            .O(N__41579),
            .I(N__41564));
    LocalMux I__9417 (
            .O(N__41576),
            .I(N__41557));
    LocalMux I__9416 (
            .O(N__41573),
            .I(N__41557));
    LocalMux I__9415 (
            .O(N__41570),
            .I(N__41557));
    LocalMux I__9414 (
            .O(N__41567),
            .I(N__41554));
    LocalMux I__9413 (
            .O(N__41564),
            .I(N__41549));
    Span4Mux_v I__9412 (
            .O(N__41557),
            .I(N__41549));
    Span4Mux_h I__9411 (
            .O(N__41554),
            .I(N__41546));
    Odrv4 I__9410 (
            .O(N__41549),
            .I(measured_delay_hc_14));
    Odrv4 I__9409 (
            .O(N__41546),
            .I(measured_delay_hc_14));
    CascadeMux I__9408 (
            .O(N__41541),
            .I(N__41535));
    CascadeMux I__9407 (
            .O(N__41540),
            .I(N__41532));
    CascadeMux I__9406 (
            .O(N__41539),
            .I(N__41529));
    CascadeMux I__9405 (
            .O(N__41538),
            .I(N__41526));
    InMux I__9404 (
            .O(N__41535),
            .I(N__41518));
    InMux I__9403 (
            .O(N__41532),
            .I(N__41501));
    InMux I__9402 (
            .O(N__41529),
            .I(N__41501));
    InMux I__9401 (
            .O(N__41526),
            .I(N__41501));
    InMux I__9400 (
            .O(N__41525),
            .I(N__41501));
    InMux I__9399 (
            .O(N__41524),
            .I(N__41501));
    InMux I__9398 (
            .O(N__41523),
            .I(N__41501));
    InMux I__9397 (
            .O(N__41522),
            .I(N__41501));
    InMux I__9396 (
            .O(N__41521),
            .I(N__41501));
    LocalMux I__9395 (
            .O(N__41518),
            .I(N__41489));
    LocalMux I__9394 (
            .O(N__41501),
            .I(N__41486));
    CascadeMux I__9393 (
            .O(N__41500),
            .I(N__41483));
    CascadeMux I__9392 (
            .O(N__41499),
            .I(N__41480));
    CascadeMux I__9391 (
            .O(N__41498),
            .I(N__41477));
    CascadeMux I__9390 (
            .O(N__41497),
            .I(N__41472));
    CascadeMux I__9389 (
            .O(N__41496),
            .I(N__41469));
    CascadeMux I__9388 (
            .O(N__41495),
            .I(N__41466));
    InMux I__9387 (
            .O(N__41494),
            .I(N__41452));
    InMux I__9386 (
            .O(N__41493),
            .I(N__41447));
    InMux I__9385 (
            .O(N__41492),
            .I(N__41447));
    Span4Mux_v I__9384 (
            .O(N__41489),
            .I(N__41442));
    Span4Mux_h I__9383 (
            .O(N__41486),
            .I(N__41442));
    InMux I__9382 (
            .O(N__41483),
            .I(N__41439));
    InMux I__9381 (
            .O(N__41480),
            .I(N__41430));
    InMux I__9380 (
            .O(N__41477),
            .I(N__41430));
    InMux I__9379 (
            .O(N__41476),
            .I(N__41430));
    InMux I__9378 (
            .O(N__41475),
            .I(N__41430));
    InMux I__9377 (
            .O(N__41472),
            .I(N__41417));
    InMux I__9376 (
            .O(N__41469),
            .I(N__41417));
    InMux I__9375 (
            .O(N__41466),
            .I(N__41417));
    InMux I__9374 (
            .O(N__41465),
            .I(N__41417));
    InMux I__9373 (
            .O(N__41464),
            .I(N__41417));
    InMux I__9372 (
            .O(N__41463),
            .I(N__41417));
    InMux I__9371 (
            .O(N__41462),
            .I(N__41412));
    InMux I__9370 (
            .O(N__41461),
            .I(N__41412));
    InMux I__9369 (
            .O(N__41460),
            .I(N__41399));
    InMux I__9368 (
            .O(N__41459),
            .I(N__41399));
    InMux I__9367 (
            .O(N__41458),
            .I(N__41399));
    InMux I__9366 (
            .O(N__41457),
            .I(N__41399));
    InMux I__9365 (
            .O(N__41456),
            .I(N__41399));
    InMux I__9364 (
            .O(N__41455),
            .I(N__41399));
    LocalMux I__9363 (
            .O(N__41452),
            .I(N__41396));
    LocalMux I__9362 (
            .O(N__41447),
            .I(N__41391));
    Span4Mux_h I__9361 (
            .O(N__41442),
            .I(N__41391));
    LocalMux I__9360 (
            .O(N__41439),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    LocalMux I__9359 (
            .O(N__41430),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    LocalMux I__9358 (
            .O(N__41417),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    LocalMux I__9357 (
            .O(N__41412),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    LocalMux I__9356 (
            .O(N__41399),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    Odrv4 I__9355 (
            .O(N__41396),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    Odrv4 I__9354 (
            .O(N__41391),
            .I(\phase_controller_inst1.stoper_hc.N_405 ));
    CascadeMux I__9353 (
            .O(N__41376),
            .I(N__41370));
    InMux I__9352 (
            .O(N__41375),
            .I(N__41367));
    InMux I__9351 (
            .O(N__41374),
            .I(N__41364));
    InMux I__9350 (
            .O(N__41373),
            .I(N__41361));
    InMux I__9349 (
            .O(N__41370),
            .I(N__41357));
    LocalMux I__9348 (
            .O(N__41367),
            .I(N__41354));
    LocalMux I__9347 (
            .O(N__41364),
            .I(N__41349));
    LocalMux I__9346 (
            .O(N__41361),
            .I(N__41349));
    InMux I__9345 (
            .O(N__41360),
            .I(N__41346));
    LocalMux I__9344 (
            .O(N__41357),
            .I(N__41343));
    Span4Mux_h I__9343 (
            .O(N__41354),
            .I(N__41340));
    Span12Mux_s11_h I__9342 (
            .O(N__41349),
            .I(N__41337));
    LocalMux I__9341 (
            .O(N__41346),
            .I(measured_delay_hc_9));
    Odrv4 I__9340 (
            .O(N__41343),
            .I(measured_delay_hc_9));
    Odrv4 I__9339 (
            .O(N__41340),
            .I(measured_delay_hc_9));
    Odrv12 I__9338 (
            .O(N__41337),
            .I(measured_delay_hc_9));
    CascadeMux I__9337 (
            .O(N__41328),
            .I(N__41325));
    InMux I__9336 (
            .O(N__41325),
            .I(N__41322));
    LocalMux I__9335 (
            .O(N__41322),
            .I(N__41318));
    InMux I__9334 (
            .O(N__41321),
            .I(N__41315));
    Span4Mux_h I__9333 (
            .O(N__41318),
            .I(N__41312));
    LocalMux I__9332 (
            .O(N__41315),
            .I(N__41307));
    Span4Mux_v I__9331 (
            .O(N__41312),
            .I(N__41307));
    Odrv4 I__9330 (
            .O(N__41307),
            .I(measured_delay_hc_30));
    InMux I__9329 (
            .O(N__41304),
            .I(N__41301));
    LocalMux I__9328 (
            .O(N__41301),
            .I(N__41298));
    Odrv4 I__9327 (
            .O(N__41298),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6Z0Z_19 ));
    CascadeMux I__9326 (
            .O(N__41295),
            .I(N__41289));
    InMux I__9325 (
            .O(N__41294),
            .I(N__41286));
    InMux I__9324 (
            .O(N__41293),
            .I(N__41283));
    CascadeMux I__9323 (
            .O(N__41292),
            .I(N__41279));
    InMux I__9322 (
            .O(N__41289),
            .I(N__41276));
    LocalMux I__9321 (
            .O(N__41286),
            .I(N__41271));
    LocalMux I__9320 (
            .O(N__41283),
            .I(N__41271));
    InMux I__9319 (
            .O(N__41282),
            .I(N__41268));
    InMux I__9318 (
            .O(N__41279),
            .I(N__41265));
    LocalMux I__9317 (
            .O(N__41276),
            .I(N__41258));
    Span4Mux_v I__9316 (
            .O(N__41271),
            .I(N__41258));
    LocalMux I__9315 (
            .O(N__41268),
            .I(N__41258));
    LocalMux I__9314 (
            .O(N__41265),
            .I(measured_delay_hc_6));
    Odrv4 I__9313 (
            .O(N__41258),
            .I(measured_delay_hc_6));
    InMux I__9312 (
            .O(N__41253),
            .I(N__41249));
    InMux I__9311 (
            .O(N__41252),
            .I(N__41246));
    LocalMux I__9310 (
            .O(N__41249),
            .I(measured_delay_hc_29));
    LocalMux I__9309 (
            .O(N__41246),
            .I(measured_delay_hc_29));
    InMux I__9308 (
            .O(N__41241),
            .I(N__41235));
    InMux I__9307 (
            .O(N__41240),
            .I(N__41232));
    InMux I__9306 (
            .O(N__41239),
            .I(N__41229));
    CascadeMux I__9305 (
            .O(N__41238),
            .I(N__41226));
    LocalMux I__9304 (
            .O(N__41235),
            .I(N__41219));
    LocalMux I__9303 (
            .O(N__41232),
            .I(N__41219));
    LocalMux I__9302 (
            .O(N__41229),
            .I(N__41216));
    InMux I__9301 (
            .O(N__41226),
            .I(N__41213));
    InMux I__9300 (
            .O(N__41225),
            .I(N__41208));
    InMux I__9299 (
            .O(N__41224),
            .I(N__41208));
    Span4Mux_v I__9298 (
            .O(N__41219),
            .I(N__41203));
    Span4Mux_v I__9297 (
            .O(N__41216),
            .I(N__41203));
    LocalMux I__9296 (
            .O(N__41213),
            .I(measured_delay_hc_7));
    LocalMux I__9295 (
            .O(N__41208),
            .I(measured_delay_hc_7));
    Odrv4 I__9294 (
            .O(N__41203),
            .I(measured_delay_hc_7));
    InMux I__9293 (
            .O(N__41196),
            .I(N__41192));
    InMux I__9292 (
            .O(N__41195),
            .I(N__41188));
    LocalMux I__9291 (
            .O(N__41192),
            .I(N__41183));
    InMux I__9290 (
            .O(N__41191),
            .I(N__41180));
    LocalMux I__9289 (
            .O(N__41188),
            .I(N__41177));
    CascadeMux I__9288 (
            .O(N__41187),
            .I(N__41174));
    InMux I__9287 (
            .O(N__41186),
            .I(N__41171));
    Span4Mux_h I__9286 (
            .O(N__41183),
            .I(N__41168));
    LocalMux I__9285 (
            .O(N__41180),
            .I(N__41163));
    Span4Mux_v I__9284 (
            .O(N__41177),
            .I(N__41163));
    InMux I__9283 (
            .O(N__41174),
            .I(N__41160));
    LocalMux I__9282 (
            .O(N__41171),
            .I(measured_delay_hc_5));
    Odrv4 I__9281 (
            .O(N__41168),
            .I(measured_delay_hc_5));
    Odrv4 I__9280 (
            .O(N__41163),
            .I(measured_delay_hc_5));
    LocalMux I__9279 (
            .O(N__41160),
            .I(measured_delay_hc_5));
    InMux I__9278 (
            .O(N__41151),
            .I(N__41148));
    LocalMux I__9277 (
            .O(N__41148),
            .I(N__41145));
    Odrv4 I__9276 (
            .O(N__41145),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3Z0Z_18 ));
    CascadeMux I__9275 (
            .O(N__41142),
            .I(N__41139));
    InMux I__9274 (
            .O(N__41139),
            .I(N__41136));
    LocalMux I__9273 (
            .O(N__41136),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3Z0Z_2 ));
    InMux I__9272 (
            .O(N__41133),
            .I(N__41130));
    LocalMux I__9271 (
            .O(N__41130),
            .I(\phase_controller_inst1.stoper_hc.N_388 ));
    CascadeMux I__9270 (
            .O(N__41127),
            .I(\phase_controller_inst1.stoper_hc.N_405_cascade_ ));
    InMux I__9269 (
            .O(N__41124),
            .I(N__41120));
    InMux I__9268 (
            .O(N__41123),
            .I(N__41115));
    LocalMux I__9267 (
            .O(N__41120),
            .I(N__41112));
    InMux I__9266 (
            .O(N__41119),
            .I(N__41109));
    InMux I__9265 (
            .O(N__41118),
            .I(N__41106));
    LocalMux I__9264 (
            .O(N__41115),
            .I(N__41103));
    Span4Mux_h I__9263 (
            .O(N__41112),
            .I(N__41098));
    LocalMux I__9262 (
            .O(N__41109),
            .I(N__41098));
    LocalMux I__9261 (
            .O(N__41106),
            .I(N__41092));
    Span4Mux_v I__9260 (
            .O(N__41103),
            .I(N__41092));
    Span4Mux_v I__9259 (
            .O(N__41098),
            .I(N__41089));
    InMux I__9258 (
            .O(N__41097),
            .I(N__41086));
    Odrv4 I__9257 (
            .O(N__41092),
            .I(measured_delay_hc_4));
    Odrv4 I__9256 (
            .O(N__41089),
            .I(measured_delay_hc_4));
    LocalMux I__9255 (
            .O(N__41086),
            .I(measured_delay_hc_4));
    CascadeMux I__9254 (
            .O(N__41079),
            .I(N__41076));
    InMux I__9253 (
            .O(N__41076),
            .I(N__41072));
    CascadeMux I__9252 (
            .O(N__41075),
            .I(N__41066));
    LocalMux I__9251 (
            .O(N__41072),
            .I(N__41063));
    InMux I__9250 (
            .O(N__41071),
            .I(N__41060));
    InMux I__9249 (
            .O(N__41070),
            .I(N__41057));
    InMux I__9248 (
            .O(N__41069),
            .I(N__41054));
    InMux I__9247 (
            .O(N__41066),
            .I(N__41051));
    Span4Mux_v I__9246 (
            .O(N__41063),
            .I(N__41046));
    LocalMux I__9245 (
            .O(N__41060),
            .I(N__41046));
    LocalMux I__9244 (
            .O(N__41057),
            .I(N__41041));
    LocalMux I__9243 (
            .O(N__41054),
            .I(N__41041));
    LocalMux I__9242 (
            .O(N__41051),
            .I(measured_delay_hc_10));
    Odrv4 I__9241 (
            .O(N__41046),
            .I(measured_delay_hc_10));
    Odrv4 I__9240 (
            .O(N__41041),
            .I(measured_delay_hc_10));
    InMux I__9239 (
            .O(N__41034),
            .I(N__41031));
    LocalMux I__9238 (
            .O(N__41031),
            .I(N__41025));
    CascadeMux I__9237 (
            .O(N__41030),
            .I(N__41022));
    CascadeMux I__9236 (
            .O(N__41029),
            .I(N__41019));
    InMux I__9235 (
            .O(N__41028),
            .I(N__41015));
    Span4Mux_h I__9234 (
            .O(N__41025),
            .I(N__41012));
    InMux I__9233 (
            .O(N__41022),
            .I(N__41009));
    InMux I__9232 (
            .O(N__41019),
            .I(N__41004));
    InMux I__9231 (
            .O(N__41018),
            .I(N__41004));
    LocalMux I__9230 (
            .O(N__41015),
            .I(N__41001));
    Odrv4 I__9229 (
            .O(N__41012),
            .I(measured_delay_hc_11));
    LocalMux I__9228 (
            .O(N__41009),
            .I(measured_delay_hc_11));
    LocalMux I__9227 (
            .O(N__41004),
            .I(measured_delay_hc_11));
    Odrv4 I__9226 (
            .O(N__41001),
            .I(measured_delay_hc_11));
    CascadeMux I__9225 (
            .O(N__40992),
            .I(N__40987));
    InMux I__9224 (
            .O(N__40991),
            .I(N__40984));
    CascadeMux I__9223 (
            .O(N__40990),
            .I(N__40981));
    InMux I__9222 (
            .O(N__40987),
            .I(N__40978));
    LocalMux I__9221 (
            .O(N__40984),
            .I(N__40975));
    InMux I__9220 (
            .O(N__40981),
            .I(N__40972));
    LocalMux I__9219 (
            .O(N__40978),
            .I(N__40967));
    Span4Mux_h I__9218 (
            .O(N__40975),
            .I(N__40962));
    LocalMux I__9217 (
            .O(N__40972),
            .I(N__40962));
    InMux I__9216 (
            .O(N__40971),
            .I(N__40957));
    InMux I__9215 (
            .O(N__40970),
            .I(N__40957));
    Odrv4 I__9214 (
            .O(N__40967),
            .I(measured_delay_hc_12));
    Odrv4 I__9213 (
            .O(N__40962),
            .I(measured_delay_hc_12));
    LocalMux I__9212 (
            .O(N__40957),
            .I(measured_delay_hc_12));
    InMux I__9211 (
            .O(N__40950),
            .I(N__40947));
    LocalMux I__9210 (
            .O(N__40947),
            .I(N__40942));
    InMux I__9209 (
            .O(N__40946),
            .I(N__40939));
    InMux I__9208 (
            .O(N__40945),
            .I(N__40934));
    Span4Mux_h I__9207 (
            .O(N__40942),
            .I(N__40929));
    LocalMux I__9206 (
            .O(N__40939),
            .I(N__40929));
    InMux I__9205 (
            .O(N__40938),
            .I(N__40926));
    CascadeMux I__9204 (
            .O(N__40937),
            .I(N__40923));
    LocalMux I__9203 (
            .O(N__40934),
            .I(N__40918));
    Span4Mux_h I__9202 (
            .O(N__40929),
            .I(N__40918));
    LocalMux I__9201 (
            .O(N__40926),
            .I(N__40915));
    InMux I__9200 (
            .O(N__40923),
            .I(N__40912));
    Span4Mux_v I__9199 (
            .O(N__40918),
            .I(N__40907));
    Span4Mux_h I__9198 (
            .O(N__40915),
            .I(N__40907));
    LocalMux I__9197 (
            .O(N__40912),
            .I(measured_delay_hc_8));
    Odrv4 I__9196 (
            .O(N__40907),
            .I(measured_delay_hc_8));
    InMux I__9195 (
            .O(N__40902),
            .I(N__40899));
    LocalMux I__9194 (
            .O(N__40899),
            .I(N__40895));
    InMux I__9193 (
            .O(N__40898),
            .I(N__40892));
    Span4Mux_h I__9192 (
            .O(N__40895),
            .I(N__40889));
    LocalMux I__9191 (
            .O(N__40892),
            .I(N__40886));
    Odrv4 I__9190 (
            .O(N__40889),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1 ));
    Odrv4 I__9189 (
            .O(N__40886),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1 ));
    CascadeMux I__9188 (
            .O(N__40881),
            .I(N__40878));
    InMux I__9187 (
            .O(N__40878),
            .I(N__40875));
    LocalMux I__9186 (
            .O(N__40875),
            .I(N__40872));
    Span4Mux_h I__9185 (
            .O(N__40872),
            .I(N__40869));
    Odrv4 I__9184 (
            .O(N__40869),
            .I(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ));
    InMux I__9183 (
            .O(N__40866),
            .I(N__40862));
    InMux I__9182 (
            .O(N__40865),
            .I(N__40859));
    LocalMux I__9181 (
            .O(N__40862),
            .I(N__40855));
    LocalMux I__9180 (
            .O(N__40859),
            .I(N__40852));
    InMux I__9179 (
            .O(N__40858),
            .I(N__40849));
    Odrv4 I__9178 (
            .O(N__40855),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    Odrv4 I__9177 (
            .O(N__40852),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    LocalMux I__9176 (
            .O(N__40849),
            .I(\delay_measurement_inst.hc_stateZ0Z_0 ));
    InMux I__9175 (
            .O(N__40842),
            .I(N__40839));
    LocalMux I__9174 (
            .O(N__40839),
            .I(N__40834));
    InMux I__9173 (
            .O(N__40838),
            .I(N__40831));
    InMux I__9172 (
            .O(N__40837),
            .I(N__40828));
    Span4Mux_h I__9171 (
            .O(N__40834),
            .I(N__40825));
    LocalMux I__9170 (
            .O(N__40831),
            .I(N__40822));
    LocalMux I__9169 (
            .O(N__40828),
            .I(N__40819));
    Sp12to4 I__9168 (
            .O(N__40825),
            .I(N__40816));
    Sp12to4 I__9167 (
            .O(N__40822),
            .I(N__40813));
    Span4Mux_h I__9166 (
            .O(N__40819),
            .I(N__40810));
    Span12Mux_v I__9165 (
            .O(N__40816),
            .I(N__40807));
    Span12Mux_s10_v I__9164 (
            .O(N__40813),
            .I(N__40804));
    Odrv4 I__9163 (
            .O(N__40810),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv12 I__9162 (
            .O(N__40807),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv12 I__9161 (
            .O(N__40804),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CascadeMux I__9160 (
            .O(N__40797),
            .I(\phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa_cascade_ ));
    InMux I__9159 (
            .O(N__40794),
            .I(N__40789));
    InMux I__9158 (
            .O(N__40793),
            .I(N__40786));
    InMux I__9157 (
            .O(N__40792),
            .I(N__40783));
    LocalMux I__9156 (
            .O(N__40789),
            .I(N__40777));
    LocalMux I__9155 (
            .O(N__40786),
            .I(N__40777));
    LocalMux I__9154 (
            .O(N__40783),
            .I(N__40774));
    InMux I__9153 (
            .O(N__40782),
            .I(N__40771));
    Span12Mux_h I__9152 (
            .O(N__40777),
            .I(N__40768));
    Odrv12 I__9151 (
            .O(N__40774),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__9150 (
            .O(N__40771),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__9149 (
            .O(N__40768),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__9148 (
            .O(N__40761),
            .I(N__40756));
    InMux I__9147 (
            .O(N__40760),
            .I(N__40753));
    InMux I__9146 (
            .O(N__40759),
            .I(N__40750));
    LocalMux I__9145 (
            .O(N__40756),
            .I(N__40744));
    LocalMux I__9144 (
            .O(N__40753),
            .I(N__40744));
    LocalMux I__9143 (
            .O(N__40750),
            .I(N__40741));
    InMux I__9142 (
            .O(N__40749),
            .I(N__40738));
    Span4Mux_v I__9141 (
            .O(N__40744),
            .I(N__40733));
    Span4Mux_h I__9140 (
            .O(N__40741),
            .I(N__40733));
    LocalMux I__9139 (
            .O(N__40738),
            .I(N__40730));
    Span4Mux_v I__9138 (
            .O(N__40733),
            .I(N__40727));
    Span4Mux_v I__9137 (
            .O(N__40730),
            .I(N__40724));
    Odrv4 I__9136 (
            .O(N__40727),
            .I(delay_hc_d2));
    Odrv4 I__9135 (
            .O(N__40724),
            .I(delay_hc_d2));
    InMux I__9134 (
            .O(N__40719),
            .I(N__40716));
    LocalMux I__9133 (
            .O(N__40716),
            .I(N__40712));
    InMux I__9132 (
            .O(N__40715),
            .I(N__40709));
    Span12Mux_h I__9131 (
            .O(N__40712),
            .I(N__40705));
    LocalMux I__9130 (
            .O(N__40709),
            .I(N__40702));
    InMux I__9129 (
            .O(N__40708),
            .I(N__40699));
    Odrv12 I__9128 (
            .O(N__40705),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    Odrv4 I__9127 (
            .O(N__40702),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    LocalMux I__9126 (
            .O(N__40699),
            .I(\delay_measurement_inst.prev_hc_sigZ0 ));
    CascadeMux I__9125 (
            .O(N__40692),
            .I(N__40688));
    CascadeMux I__9124 (
            .O(N__40691),
            .I(N__40685));
    InMux I__9123 (
            .O(N__40688),
            .I(N__40679));
    InMux I__9122 (
            .O(N__40685),
            .I(N__40679));
    InMux I__9121 (
            .O(N__40684),
            .I(N__40676));
    LocalMux I__9120 (
            .O(N__40679),
            .I(N__40673));
    LocalMux I__9119 (
            .O(N__40676),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__9118 (
            .O(N__40673),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__9117 (
            .O(N__40668),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9116 (
            .O(N__40665),
            .I(N__40661));
    CascadeMux I__9115 (
            .O(N__40664),
            .I(N__40658));
    LocalMux I__9114 (
            .O(N__40661),
            .I(N__40654));
    InMux I__9113 (
            .O(N__40658),
            .I(N__40651));
    InMux I__9112 (
            .O(N__40657),
            .I(N__40648));
    Span4Mux_v I__9111 (
            .O(N__40654),
            .I(N__40643));
    LocalMux I__9110 (
            .O(N__40651),
            .I(N__40643));
    LocalMux I__9109 (
            .O(N__40648),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__9108 (
            .O(N__40643),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__9107 (
            .O(N__40638),
            .I(bfn_17_11_0_));
    CascadeMux I__9106 (
            .O(N__40635),
            .I(N__40632));
    InMux I__9105 (
            .O(N__40632),
            .I(N__40629));
    LocalMux I__9104 (
            .O(N__40629),
            .I(N__40624));
    InMux I__9103 (
            .O(N__40628),
            .I(N__40621));
    InMux I__9102 (
            .O(N__40627),
            .I(N__40618));
    Span4Mux_v I__9101 (
            .O(N__40624),
            .I(N__40615));
    LocalMux I__9100 (
            .O(N__40621),
            .I(N__40612));
    LocalMux I__9099 (
            .O(N__40618),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__9098 (
            .O(N__40615),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__9097 (
            .O(N__40612),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__9096 (
            .O(N__40605),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__9095 (
            .O(N__40602),
            .I(N__40598));
    CascadeMux I__9094 (
            .O(N__40601),
            .I(N__40595));
    InMux I__9093 (
            .O(N__40598),
            .I(N__40589));
    InMux I__9092 (
            .O(N__40595),
            .I(N__40589));
    InMux I__9091 (
            .O(N__40594),
            .I(N__40586));
    LocalMux I__9090 (
            .O(N__40589),
            .I(N__40583));
    LocalMux I__9089 (
            .O(N__40586),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv4 I__9088 (
            .O(N__40583),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__9087 (
            .O(N__40578),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__9086 (
            .O(N__40575),
            .I(N__40568));
    InMux I__9085 (
            .O(N__40574),
            .I(N__40568));
    InMux I__9084 (
            .O(N__40573),
            .I(N__40565));
    LocalMux I__9083 (
            .O(N__40568),
            .I(N__40562));
    LocalMux I__9082 (
            .O(N__40565),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__9081 (
            .O(N__40562),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__9080 (
            .O(N__40557),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9079 (
            .O(N__40554),
            .I(N__40551));
    LocalMux I__9078 (
            .O(N__40551),
            .I(N__40547));
    InMux I__9077 (
            .O(N__40550),
            .I(N__40544));
    Span4Mux_h I__9076 (
            .O(N__40547),
            .I(N__40541));
    LocalMux I__9075 (
            .O(N__40544),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv4 I__9074 (
            .O(N__40541),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__9073 (
            .O(N__40536),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__9072 (
            .O(N__40533),
            .I(N__40513));
    InMux I__9071 (
            .O(N__40532),
            .I(N__40513));
    InMux I__9070 (
            .O(N__40531),
            .I(N__40513));
    InMux I__9069 (
            .O(N__40530),
            .I(N__40513));
    InMux I__9068 (
            .O(N__40529),
            .I(N__40504));
    InMux I__9067 (
            .O(N__40528),
            .I(N__40504));
    InMux I__9066 (
            .O(N__40527),
            .I(N__40504));
    InMux I__9065 (
            .O(N__40526),
            .I(N__40504));
    InMux I__9064 (
            .O(N__40525),
            .I(N__40495));
    InMux I__9063 (
            .O(N__40524),
            .I(N__40495));
    InMux I__9062 (
            .O(N__40523),
            .I(N__40495));
    InMux I__9061 (
            .O(N__40522),
            .I(N__40495));
    LocalMux I__9060 (
            .O(N__40513),
            .I(N__40478));
    LocalMux I__9059 (
            .O(N__40504),
            .I(N__40478));
    LocalMux I__9058 (
            .O(N__40495),
            .I(N__40478));
    InMux I__9057 (
            .O(N__40494),
            .I(N__40473));
    InMux I__9056 (
            .O(N__40493),
            .I(N__40473));
    InMux I__9055 (
            .O(N__40492),
            .I(N__40464));
    InMux I__9054 (
            .O(N__40491),
            .I(N__40464));
    InMux I__9053 (
            .O(N__40490),
            .I(N__40464));
    InMux I__9052 (
            .O(N__40489),
            .I(N__40464));
    InMux I__9051 (
            .O(N__40488),
            .I(N__40447));
    InMux I__9050 (
            .O(N__40487),
            .I(N__40447));
    InMux I__9049 (
            .O(N__40486),
            .I(N__40447));
    InMux I__9048 (
            .O(N__40485),
            .I(N__40447));
    Span4Mux_v I__9047 (
            .O(N__40478),
            .I(N__40440));
    LocalMux I__9046 (
            .O(N__40473),
            .I(N__40440));
    LocalMux I__9045 (
            .O(N__40464),
            .I(N__40440));
    InMux I__9044 (
            .O(N__40463),
            .I(N__40431));
    InMux I__9043 (
            .O(N__40462),
            .I(N__40431));
    InMux I__9042 (
            .O(N__40461),
            .I(N__40431));
    InMux I__9041 (
            .O(N__40460),
            .I(N__40431));
    InMux I__9040 (
            .O(N__40459),
            .I(N__40422));
    InMux I__9039 (
            .O(N__40458),
            .I(N__40422));
    InMux I__9038 (
            .O(N__40457),
            .I(N__40422));
    InMux I__9037 (
            .O(N__40456),
            .I(N__40422));
    LocalMux I__9036 (
            .O(N__40447),
            .I(N__40417));
    Span4Mux_v I__9035 (
            .O(N__40440),
            .I(N__40417));
    LocalMux I__9034 (
            .O(N__40431),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    LocalMux I__9033 (
            .O(N__40422),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9032 (
            .O(N__40417),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9031 (
            .O(N__40410),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CascadeMux I__9030 (
            .O(N__40407),
            .I(N__40404));
    InMux I__9029 (
            .O(N__40404),
            .I(N__40401));
    LocalMux I__9028 (
            .O(N__40401),
            .I(N__40397));
    InMux I__9027 (
            .O(N__40400),
            .I(N__40394));
    Span4Mux_h I__9026 (
            .O(N__40397),
            .I(N__40391));
    LocalMux I__9025 (
            .O(N__40394),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv4 I__9024 (
            .O(N__40391),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__9023 (
            .O(N__40386),
            .I(N__40382));
    CEMux I__9022 (
            .O(N__40385),
            .I(N__40379));
    LocalMux I__9021 (
            .O(N__40382),
            .I(N__40372));
    LocalMux I__9020 (
            .O(N__40379),
            .I(N__40372));
    CEMux I__9019 (
            .O(N__40378),
            .I(N__40369));
    CEMux I__9018 (
            .O(N__40377),
            .I(N__40366));
    Span4Mux_v I__9017 (
            .O(N__40372),
            .I(N__40363));
    LocalMux I__9016 (
            .O(N__40369),
            .I(N__40358));
    LocalMux I__9015 (
            .O(N__40366),
            .I(N__40358));
    Span4Mux_h I__9014 (
            .O(N__40363),
            .I(N__40353));
    Span4Mux_v I__9013 (
            .O(N__40358),
            .I(N__40353));
    Span4Mux_h I__9012 (
            .O(N__40353),
            .I(N__40350));
    Odrv4 I__9011 (
            .O(N__40350),
            .I(\delay_measurement_inst.delay_tr_timer.N_464_i ));
    InMux I__9010 (
            .O(N__40347),
            .I(N__40344));
    LocalMux I__9009 (
            .O(N__40344),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9008 (
            .O(N__40341),
            .I(N__40338));
    LocalMux I__9007 (
            .O(N__40338),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__9006 (
            .O(N__40335),
            .I(N__40332));
    LocalMux I__9005 (
            .O(N__40332),
            .I(N__40329));
    Odrv4 I__9004 (
            .O(N__40329),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ));
    CascadeMux I__9003 (
            .O(N__40326),
            .I(N__40322));
    CascadeMux I__9002 (
            .O(N__40325),
            .I(N__40319));
    InMux I__9001 (
            .O(N__40322),
            .I(N__40314));
    InMux I__9000 (
            .O(N__40319),
            .I(N__40314));
    LocalMux I__8999 (
            .O(N__40314),
            .I(N__40310));
    InMux I__8998 (
            .O(N__40313),
            .I(N__40307));
    Span4Mux_h I__8997 (
            .O(N__40310),
            .I(N__40304));
    LocalMux I__8996 (
            .O(N__40307),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__8995 (
            .O(N__40304),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__8994 (
            .O(N__40299),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__8993 (
            .O(N__40296),
            .I(N__40292));
    CascadeMux I__8992 (
            .O(N__40295),
            .I(N__40289));
    InMux I__8991 (
            .O(N__40292),
            .I(N__40283));
    InMux I__8990 (
            .O(N__40289),
            .I(N__40283));
    InMux I__8989 (
            .O(N__40288),
            .I(N__40280));
    LocalMux I__8988 (
            .O(N__40283),
            .I(N__40277));
    LocalMux I__8987 (
            .O(N__40280),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__8986 (
            .O(N__40277),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__8985 (
            .O(N__40272),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__8984 (
            .O(N__40269),
            .I(N__40265));
    InMux I__8983 (
            .O(N__40268),
            .I(N__40262));
    LocalMux I__8982 (
            .O(N__40265),
            .I(N__40259));
    LocalMux I__8981 (
            .O(N__40262),
            .I(N__40255));
    Span4Mux_v I__8980 (
            .O(N__40259),
            .I(N__40252));
    InMux I__8979 (
            .O(N__40258),
            .I(N__40249));
    Span4Mux_h I__8978 (
            .O(N__40255),
            .I(N__40246));
    Odrv4 I__8977 (
            .O(N__40252),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__8976 (
            .O(N__40249),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__8975 (
            .O(N__40246),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__8974 (
            .O(N__40239),
            .I(bfn_17_10_0_));
    InMux I__8973 (
            .O(N__40236),
            .I(N__40233));
    LocalMux I__8972 (
            .O(N__40233),
            .I(N__40228));
    InMux I__8971 (
            .O(N__40232),
            .I(N__40225));
    InMux I__8970 (
            .O(N__40231),
            .I(N__40222));
    Span4Mux_v I__8969 (
            .O(N__40228),
            .I(N__40217));
    LocalMux I__8968 (
            .O(N__40225),
            .I(N__40217));
    LocalMux I__8967 (
            .O(N__40222),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__8966 (
            .O(N__40217),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__8965 (
            .O(N__40212),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__8964 (
            .O(N__40209),
            .I(N__40205));
    CascadeMux I__8963 (
            .O(N__40208),
            .I(N__40202));
    InMux I__8962 (
            .O(N__40205),
            .I(N__40196));
    InMux I__8961 (
            .O(N__40202),
            .I(N__40196));
    InMux I__8960 (
            .O(N__40201),
            .I(N__40193));
    LocalMux I__8959 (
            .O(N__40196),
            .I(N__40190));
    LocalMux I__8958 (
            .O(N__40193),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv4 I__8957 (
            .O(N__40190),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__8956 (
            .O(N__40185),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__8955 (
            .O(N__40182),
            .I(N__40178));
    CascadeMux I__8954 (
            .O(N__40181),
            .I(N__40175));
    InMux I__8953 (
            .O(N__40178),
            .I(N__40170));
    InMux I__8952 (
            .O(N__40175),
            .I(N__40170));
    LocalMux I__8951 (
            .O(N__40170),
            .I(N__40166));
    InMux I__8950 (
            .O(N__40169),
            .I(N__40163));
    Span4Mux_h I__8949 (
            .O(N__40166),
            .I(N__40160));
    LocalMux I__8948 (
            .O(N__40163),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__8947 (
            .O(N__40160),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__8946 (
            .O(N__40155),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__8945 (
            .O(N__40152),
            .I(N__40148));
    InMux I__8944 (
            .O(N__40151),
            .I(N__40145));
    InMux I__8943 (
            .O(N__40148),
            .I(N__40141));
    LocalMux I__8942 (
            .O(N__40145),
            .I(N__40138));
    InMux I__8941 (
            .O(N__40144),
            .I(N__40135));
    LocalMux I__8940 (
            .O(N__40141),
            .I(N__40130));
    Span4Mux_h I__8939 (
            .O(N__40138),
            .I(N__40130));
    LocalMux I__8938 (
            .O(N__40135),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__8937 (
            .O(N__40130),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__8936 (
            .O(N__40125),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__8935 (
            .O(N__40122),
            .I(N__40115));
    InMux I__8934 (
            .O(N__40121),
            .I(N__40115));
    InMux I__8933 (
            .O(N__40120),
            .I(N__40112));
    LocalMux I__8932 (
            .O(N__40115),
            .I(N__40109));
    LocalMux I__8931 (
            .O(N__40112),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv4 I__8930 (
            .O(N__40109),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__8929 (
            .O(N__40104),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__8928 (
            .O(N__40101),
            .I(N__40094));
    InMux I__8927 (
            .O(N__40100),
            .I(N__40094));
    InMux I__8926 (
            .O(N__40099),
            .I(N__40091));
    LocalMux I__8925 (
            .O(N__40094),
            .I(N__40088));
    LocalMux I__8924 (
            .O(N__40091),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__8923 (
            .O(N__40088),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__8922 (
            .O(N__40083),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__8921 (
            .O(N__40080),
            .I(N__40073));
    InMux I__8920 (
            .O(N__40079),
            .I(N__40073));
    InMux I__8919 (
            .O(N__40078),
            .I(N__40070));
    LocalMux I__8918 (
            .O(N__40073),
            .I(N__40067));
    LocalMux I__8917 (
            .O(N__40070),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__8916 (
            .O(N__40067),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__8915 (
            .O(N__40062),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__8914 (
            .O(N__40059),
            .I(N__40055));
    CascadeMux I__8913 (
            .O(N__40058),
            .I(N__40052));
    InMux I__8912 (
            .O(N__40055),
            .I(N__40047));
    InMux I__8911 (
            .O(N__40052),
            .I(N__40047));
    LocalMux I__8910 (
            .O(N__40047),
            .I(N__40043));
    InMux I__8909 (
            .O(N__40046),
            .I(N__40040));
    Span4Mux_h I__8908 (
            .O(N__40043),
            .I(N__40037));
    LocalMux I__8907 (
            .O(N__40040),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__8906 (
            .O(N__40037),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__8905 (
            .O(N__40032),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__8904 (
            .O(N__40029),
            .I(N__40025));
    CascadeMux I__8903 (
            .O(N__40028),
            .I(N__40022));
    LocalMux I__8902 (
            .O(N__40025),
            .I(N__40018));
    InMux I__8901 (
            .O(N__40022),
            .I(N__40015));
    InMux I__8900 (
            .O(N__40021),
            .I(N__40012));
    Span4Mux_v I__8899 (
            .O(N__40018),
            .I(N__40007));
    LocalMux I__8898 (
            .O(N__40015),
            .I(N__40007));
    LocalMux I__8897 (
            .O(N__40012),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__8896 (
            .O(N__40007),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__8895 (
            .O(N__40002),
            .I(bfn_17_9_0_));
    CascadeMux I__8894 (
            .O(N__39999),
            .I(N__39996));
    InMux I__8893 (
            .O(N__39996),
            .I(N__39992));
    InMux I__8892 (
            .O(N__39995),
            .I(N__39988));
    LocalMux I__8891 (
            .O(N__39992),
            .I(N__39985));
    InMux I__8890 (
            .O(N__39991),
            .I(N__39982));
    LocalMux I__8889 (
            .O(N__39988),
            .I(N__39977));
    Span4Mux_v I__8888 (
            .O(N__39985),
            .I(N__39977));
    LocalMux I__8887 (
            .O(N__39982),
            .I(N__39974));
    Odrv4 I__8886 (
            .O(N__39977),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv4 I__8885 (
            .O(N__39974),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__8884 (
            .O(N__39969),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__8883 (
            .O(N__39966),
            .I(N__39962));
    CascadeMux I__8882 (
            .O(N__39965),
            .I(N__39959));
    InMux I__8881 (
            .O(N__39962),
            .I(N__39953));
    InMux I__8880 (
            .O(N__39959),
            .I(N__39953));
    InMux I__8879 (
            .O(N__39958),
            .I(N__39950));
    LocalMux I__8878 (
            .O(N__39953),
            .I(N__39947));
    LocalMux I__8877 (
            .O(N__39950),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__8876 (
            .O(N__39947),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__8875 (
            .O(N__39942),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__8874 (
            .O(N__39939),
            .I(N__39932));
    InMux I__8873 (
            .O(N__39938),
            .I(N__39932));
    InMux I__8872 (
            .O(N__39937),
            .I(N__39929));
    LocalMux I__8871 (
            .O(N__39932),
            .I(N__39926));
    LocalMux I__8870 (
            .O(N__39929),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__8869 (
            .O(N__39926),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__8868 (
            .O(N__39921),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__8867 (
            .O(N__39918),
            .I(N__39912));
    InMux I__8866 (
            .O(N__39917),
            .I(N__39912));
    LocalMux I__8865 (
            .O(N__39912),
            .I(N__39908));
    InMux I__8864 (
            .O(N__39911),
            .I(N__39905));
    Span4Mux_h I__8863 (
            .O(N__39908),
            .I(N__39902));
    LocalMux I__8862 (
            .O(N__39905),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv4 I__8861 (
            .O(N__39902),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__8860 (
            .O(N__39897),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__8859 (
            .O(N__39894),
            .I(N__39891));
    InMux I__8858 (
            .O(N__39891),
            .I(N__39887));
    InMux I__8857 (
            .O(N__39890),
            .I(N__39883));
    LocalMux I__8856 (
            .O(N__39887),
            .I(N__39880));
    InMux I__8855 (
            .O(N__39886),
            .I(N__39877));
    LocalMux I__8854 (
            .O(N__39883),
            .I(N__39872));
    Span4Mux_h I__8853 (
            .O(N__39880),
            .I(N__39872));
    LocalMux I__8852 (
            .O(N__39877),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv4 I__8851 (
            .O(N__39872),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__8850 (
            .O(N__39867),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__8849 (
            .O(N__39864),
            .I(N__39860));
    InMux I__8848 (
            .O(N__39863),
            .I(N__39857));
    LocalMux I__8847 (
            .O(N__39860),
            .I(N__39851));
    LocalMux I__8846 (
            .O(N__39857),
            .I(N__39851));
    InMux I__8845 (
            .O(N__39856),
            .I(N__39848));
    Sp12to4 I__8844 (
            .O(N__39851),
            .I(N__39842));
    LocalMux I__8843 (
            .O(N__39848),
            .I(N__39842));
    InMux I__8842 (
            .O(N__39847),
            .I(N__39839));
    Span12Mux_v I__8841 (
            .O(N__39842),
            .I(N__39836));
    LocalMux I__8840 (
            .O(N__39839),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__8839 (
            .O(N__39836),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    IoInMux I__8838 (
            .O(N__39831),
            .I(N__39828));
    LocalMux I__8837 (
            .O(N__39828),
            .I(N__39825));
    IoSpan4Mux I__8836 (
            .O(N__39825),
            .I(N__39822));
    IoSpan4Mux I__8835 (
            .O(N__39822),
            .I(N__39819));
    IoSpan4Mux I__8834 (
            .O(N__39819),
            .I(N__39816));
    Odrv4 I__8833 (
            .O(N__39816),
            .I(\delay_measurement_inst.delay_hc_timer.N_461_i ));
    InMux I__8832 (
            .O(N__39813),
            .I(N__39810));
    LocalMux I__8831 (
            .O(N__39810),
            .I(N__39807));
    Odrv12 I__8830 (
            .O(N__39807),
            .I(delay_hc_input_c));
    InMux I__8829 (
            .O(N__39804),
            .I(N__39801));
    LocalMux I__8828 (
            .O(N__39801),
            .I(delay_hc_d1));
    InMux I__8827 (
            .O(N__39798),
            .I(bfn_17_8_0_));
    CascadeMux I__8826 (
            .O(N__39795),
            .I(N__39792));
    InMux I__8825 (
            .O(N__39792),
            .I(N__39789));
    LocalMux I__8824 (
            .O(N__39789),
            .I(N__39785));
    InMux I__8823 (
            .O(N__39788),
            .I(N__39782));
    Span4Mux_v I__8822 (
            .O(N__39785),
            .I(N__39778));
    LocalMux I__8821 (
            .O(N__39782),
            .I(N__39775));
    InMux I__8820 (
            .O(N__39781),
            .I(N__39772));
    Span4Mux_h I__8819 (
            .O(N__39778),
            .I(N__39769));
    Odrv4 I__8818 (
            .O(N__39775),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__8817 (
            .O(N__39772),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__8816 (
            .O(N__39769),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__8815 (
            .O(N__39762),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__8814 (
            .O(N__39759),
            .I(N__39755));
    CascadeMux I__8813 (
            .O(N__39758),
            .I(N__39752));
    InMux I__8812 (
            .O(N__39755),
            .I(N__39746));
    InMux I__8811 (
            .O(N__39752),
            .I(N__39746));
    InMux I__8810 (
            .O(N__39751),
            .I(N__39743));
    LocalMux I__8809 (
            .O(N__39746),
            .I(N__39740));
    LocalMux I__8808 (
            .O(N__39743),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__8807 (
            .O(N__39740),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__8806 (
            .O(N__39735),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__8805 (
            .O(N__39732),
            .I(N__39725));
    InMux I__8804 (
            .O(N__39731),
            .I(N__39725));
    InMux I__8803 (
            .O(N__39730),
            .I(N__39722));
    LocalMux I__8802 (
            .O(N__39725),
            .I(N__39719));
    LocalMux I__8801 (
            .O(N__39722),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__8800 (
            .O(N__39719),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__8799 (
            .O(N__39714),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    CascadeMux I__8798 (
            .O(N__39711),
            .I(N__39707));
    InMux I__8797 (
            .O(N__39710),
            .I(N__39704));
    InMux I__8796 (
            .O(N__39707),
            .I(N__39700));
    LocalMux I__8795 (
            .O(N__39704),
            .I(N__39697));
    InMux I__8794 (
            .O(N__39703),
            .I(N__39694));
    LocalMux I__8793 (
            .O(N__39700),
            .I(N__39689));
    Span4Mux_h I__8792 (
            .O(N__39697),
            .I(N__39689));
    LocalMux I__8791 (
            .O(N__39694),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv4 I__8790 (
            .O(N__39689),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__8789 (
            .O(N__39684),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__8788 (
            .O(N__39681),
            .I(N__39678));
    InMux I__8787 (
            .O(N__39678),
            .I(N__39674));
    InMux I__8786 (
            .O(N__39677),
            .I(N__39670));
    LocalMux I__8785 (
            .O(N__39674),
            .I(N__39667));
    InMux I__8784 (
            .O(N__39673),
            .I(N__39664));
    LocalMux I__8783 (
            .O(N__39670),
            .I(N__39659));
    Span4Mux_h I__8782 (
            .O(N__39667),
            .I(N__39659));
    LocalMux I__8781 (
            .O(N__39664),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__8780 (
            .O(N__39659),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__8779 (
            .O(N__39654),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__8778 (
            .O(N__39651),
            .I(N__39648));
    LocalMux I__8777 (
            .O(N__39648),
            .I(N__39644));
    InMux I__8776 (
            .O(N__39647),
            .I(N__39641));
    Span4Mux_h I__8775 (
            .O(N__39644),
            .I(N__39638));
    LocalMux I__8774 (
            .O(N__39641),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__8773 (
            .O(N__39638),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__8772 (
            .O(N__39633),
            .I(N__39630));
    LocalMux I__8771 (
            .O(N__39630),
            .I(\delay_measurement_inst.delay_hc_timer.N_319 ));
    CascadeMux I__8770 (
            .O(N__39627),
            .I(\delay_measurement_inst.N_318_cascade_ ));
    InMux I__8769 (
            .O(N__39624),
            .I(N__39621));
    LocalMux I__8768 (
            .O(N__39621),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__8767 (
            .O(N__39618),
            .I(N__39615));
    LocalMux I__8766 (
            .O(N__39615),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    CascadeMux I__8765 (
            .O(N__39612),
            .I(N__39609));
    InMux I__8764 (
            .O(N__39609),
            .I(N__39606));
    LocalMux I__8763 (
            .O(N__39606),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__8762 (
            .O(N__39603),
            .I(N__39600));
    LocalMux I__8761 (
            .O(N__39600),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__8760 (
            .O(N__39597),
            .I(N__39594));
    LocalMux I__8759 (
            .O(N__39594),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_6_6 ));
    InMux I__8758 (
            .O(N__39591),
            .I(N__39588));
    LocalMux I__8757 (
            .O(N__39588),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__8756 (
            .O(N__39585),
            .I(N__39582));
    LocalMux I__8755 (
            .O(N__39582),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    CascadeMux I__8754 (
            .O(N__39579),
            .I(N__39576));
    InMux I__8753 (
            .O(N__39576),
            .I(N__39573));
    LocalMux I__8752 (
            .O(N__39573),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__8751 (
            .O(N__39570),
            .I(N__39567));
    LocalMux I__8750 (
            .O(N__39567),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__8749 (
            .O(N__39564),
            .I(N__39561));
    LocalMux I__8748 (
            .O(N__39561),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_7_6 ));
    InMux I__8747 (
            .O(N__39558),
            .I(N__39555));
    LocalMux I__8746 (
            .O(N__39555),
            .I(N__39551));
    InMux I__8745 (
            .O(N__39554),
            .I(N__39548));
    Span4Mux_h I__8744 (
            .O(N__39551),
            .I(N__39545));
    LocalMux I__8743 (
            .O(N__39548),
            .I(measured_delay_hc_21));
    Odrv4 I__8742 (
            .O(N__39545),
            .I(measured_delay_hc_21));
    InMux I__8741 (
            .O(N__39540),
            .I(N__39537));
    LocalMux I__8740 (
            .O(N__39537),
            .I(N__39534));
    Odrv4 I__8739 (
            .O(N__39534),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0Z0Z_19 ));
    InMux I__8738 (
            .O(N__39531),
            .I(N__39527));
    InMux I__8737 (
            .O(N__39530),
            .I(N__39524));
    LocalMux I__8736 (
            .O(N__39527),
            .I(N__39520));
    LocalMux I__8735 (
            .O(N__39524),
            .I(N__39517));
    InMux I__8734 (
            .O(N__39523),
            .I(N__39514));
    Span4Mux_h I__8733 (
            .O(N__39520),
            .I(N__39511));
    Odrv4 I__8732 (
            .O(N__39517),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    LocalMux I__8731 (
            .O(N__39514),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    Odrv4 I__8730 (
            .O(N__39511),
            .I(\delay_measurement_inst.elapsed_time_hc_8 ));
    CascadeMux I__8729 (
            .O(N__39504),
            .I(N__39500));
    InMux I__8728 (
            .O(N__39503),
            .I(N__39497));
    InMux I__8727 (
            .O(N__39500),
            .I(N__39494));
    LocalMux I__8726 (
            .O(N__39497),
            .I(N__39491));
    LocalMux I__8725 (
            .O(N__39494),
            .I(\delay_measurement_inst.delay_hc_timer.N_408 ));
    Odrv4 I__8724 (
            .O(N__39491),
            .I(\delay_measurement_inst.delay_hc_timer.N_408 ));
    CascadeMux I__8723 (
            .O(N__39486),
            .I(N__39483));
    InMux I__8722 (
            .O(N__39483),
            .I(N__39480));
    LocalMux I__8721 (
            .O(N__39480),
            .I(N__39476));
    InMux I__8720 (
            .O(N__39479),
            .I(N__39473));
    Span4Mux_h I__8719 (
            .O(N__39476),
            .I(N__39470));
    LocalMux I__8718 (
            .O(N__39473),
            .I(measured_delay_hc_26));
    Odrv4 I__8717 (
            .O(N__39470),
            .I(measured_delay_hc_26));
    InMux I__8716 (
            .O(N__39465),
            .I(N__39461));
    CascadeMux I__8715 (
            .O(N__39464),
            .I(N__39457));
    LocalMux I__8714 (
            .O(N__39461),
            .I(N__39454));
    InMux I__8713 (
            .O(N__39460),
            .I(N__39451));
    InMux I__8712 (
            .O(N__39457),
            .I(N__39448));
    Odrv4 I__8711 (
            .O(N__39454),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__8710 (
            .O(N__39451),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    LocalMux I__8709 (
            .O(N__39448),
            .I(\delay_measurement_inst.elapsed_time_hc_17 ));
    InMux I__8708 (
            .O(N__39441),
            .I(N__39437));
    InMux I__8707 (
            .O(N__39440),
            .I(N__39434));
    LocalMux I__8706 (
            .O(N__39437),
            .I(measured_delay_hc_20));
    LocalMux I__8705 (
            .O(N__39434),
            .I(measured_delay_hc_20));
    InMux I__8704 (
            .O(N__39429),
            .I(N__39426));
    LocalMux I__8703 (
            .O(N__39426),
            .I(N__39421));
    InMux I__8702 (
            .O(N__39425),
            .I(N__39418));
    InMux I__8701 (
            .O(N__39424),
            .I(N__39415));
    Odrv12 I__8700 (
            .O(N__39421),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__8699 (
            .O(N__39418),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    LocalMux I__8698 (
            .O(N__39415),
            .I(\delay_measurement_inst.elapsed_time_hc_4 ));
    InMux I__8697 (
            .O(N__39408),
            .I(N__39405));
    LocalMux I__8696 (
            .O(N__39405),
            .I(N__39401));
    CascadeMux I__8695 (
            .O(N__39404),
            .I(N__39398));
    Span4Mux_v I__8694 (
            .O(N__39401),
            .I(N__39394));
    InMux I__8693 (
            .O(N__39398),
            .I(N__39389));
    InMux I__8692 (
            .O(N__39397),
            .I(N__39389));
    Odrv4 I__8691 (
            .O(N__39394),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    LocalMux I__8690 (
            .O(N__39389),
            .I(\delay_measurement_inst.elapsed_time_hc_7 ));
    CascadeMux I__8689 (
            .O(N__39384),
            .I(\delay_measurement_inst.delay_hc_timer.N_318_1_cascade_ ));
    InMux I__8688 (
            .O(N__39381),
            .I(N__39378));
    LocalMux I__8687 (
            .O(N__39378),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_6 ));
    InMux I__8686 (
            .O(N__39375),
            .I(N__39372));
    LocalMux I__8685 (
            .O(N__39372),
            .I(N__39369));
    Odrv4 I__8684 (
            .O(N__39369),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_5 ));
    CascadeMux I__8683 (
            .O(N__39366),
            .I(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_9_cascade_ ));
    InMux I__8682 (
            .O(N__39363),
            .I(N__39360));
    LocalMux I__8681 (
            .O(N__39360),
            .I(\delay_measurement_inst.delay_hc_timer.N_440 ));
    InMux I__8680 (
            .O(N__39357),
            .I(N__39354));
    LocalMux I__8679 (
            .O(N__39354),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__8678 (
            .O(N__39351),
            .I(N__39348));
    LocalMux I__8677 (
            .O(N__39348),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__8676 (
            .O(N__39345),
            .I(N__39342));
    LocalMux I__8675 (
            .O(N__39342),
            .I(N__39339));
    Odrv4 I__8674 (
            .O(N__39339),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    CascadeMux I__8673 (
            .O(N__39336),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_0_6_cascade_ ));
    CascadeMux I__8672 (
            .O(N__39333),
            .I(\delay_measurement_inst.delay_hc_timer.N_328_cascade_ ));
    InMux I__8671 (
            .O(N__39330),
            .I(N__39327));
    LocalMux I__8670 (
            .O(N__39327),
            .I(N__39324));
    Odrv4 I__8669 (
            .O(N__39324),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_4 ));
    InMux I__8668 (
            .O(N__39321),
            .I(N__39318));
    LocalMux I__8667 (
            .O(N__39318),
            .I(\delay_measurement_inst.delay_hc_timer.N_318_1 ));
    InMux I__8666 (
            .O(N__39315),
            .I(N__39309));
    InMux I__8665 (
            .O(N__39314),
            .I(N__39309));
    LocalMux I__8664 (
            .O(N__39309),
            .I(N__39304));
    InMux I__8663 (
            .O(N__39308),
            .I(N__39299));
    InMux I__8662 (
            .O(N__39307),
            .I(N__39299));
    Odrv4 I__8661 (
            .O(N__39304),
            .I(\delay_measurement_inst.delay_hc_timer.N_331 ));
    LocalMux I__8660 (
            .O(N__39299),
            .I(\delay_measurement_inst.delay_hc_timer.N_331 ));
    InMux I__8659 (
            .O(N__39294),
            .I(N__39290));
    InMux I__8658 (
            .O(N__39293),
            .I(N__39287));
    LocalMux I__8657 (
            .O(N__39290),
            .I(\delay_measurement_inst.delay_hc_timer.N_328 ));
    LocalMux I__8656 (
            .O(N__39287),
            .I(\delay_measurement_inst.delay_hc_timer.N_328 ));
    InMux I__8655 (
            .O(N__39282),
            .I(N__39279));
    LocalMux I__8654 (
            .O(N__39279),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2Z0Z_18 ));
    InMux I__8653 (
            .O(N__39276),
            .I(N__39273));
    LocalMux I__8652 (
            .O(N__39273),
            .I(N__39270));
    Span4Mux_v I__8651 (
            .O(N__39270),
            .I(N__39266));
    InMux I__8650 (
            .O(N__39269),
            .I(N__39263));
    Odrv4 I__8649 (
            .O(N__39266),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    LocalMux I__8648 (
            .O(N__39263),
            .I(\delay_measurement_inst.elapsed_time_hc_12 ));
    InMux I__8647 (
            .O(N__39258),
            .I(N__39255));
    LocalMux I__8646 (
            .O(N__39255),
            .I(N__39252));
    Span4Mux_v I__8645 (
            .O(N__39252),
            .I(N__39248));
    InMux I__8644 (
            .O(N__39251),
            .I(N__39245));
    Odrv4 I__8643 (
            .O(N__39248),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    LocalMux I__8642 (
            .O(N__39245),
            .I(\delay_measurement_inst.elapsed_time_hc_11 ));
    InMux I__8641 (
            .O(N__39240),
            .I(N__39237));
    LocalMux I__8640 (
            .O(N__39237),
            .I(N__39233));
    CascadeMux I__8639 (
            .O(N__39236),
            .I(N__39230));
    Span4Mux_h I__8638 (
            .O(N__39233),
            .I(N__39227));
    InMux I__8637 (
            .O(N__39230),
            .I(N__39224));
    Odrv4 I__8636 (
            .O(N__39227),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    LocalMux I__8635 (
            .O(N__39224),
            .I(\delay_measurement_inst.elapsed_time_hc_13 ));
    InMux I__8634 (
            .O(N__39219),
            .I(N__39216));
    LocalMux I__8633 (
            .O(N__39216),
            .I(N__39212));
    InMux I__8632 (
            .O(N__39215),
            .I(N__39209));
    Odrv4 I__8631 (
            .O(N__39212),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    LocalMux I__8630 (
            .O(N__39209),
            .I(\delay_measurement_inst.elapsed_time_hc_10 ));
    InMux I__8629 (
            .O(N__39204),
            .I(N__39200));
    InMux I__8628 (
            .O(N__39203),
            .I(N__39197));
    LocalMux I__8627 (
            .O(N__39200),
            .I(N__39194));
    LocalMux I__8626 (
            .O(N__39197),
            .I(measured_delay_hc_24));
    Odrv4 I__8625 (
            .O(N__39194),
            .I(measured_delay_hc_24));
    InMux I__8624 (
            .O(N__39189),
            .I(N__39185));
    InMux I__8623 (
            .O(N__39188),
            .I(N__39182));
    LocalMux I__8622 (
            .O(N__39185),
            .I(N__39179));
    LocalMux I__8621 (
            .O(N__39182),
            .I(measured_delay_hc_23));
    Odrv12 I__8620 (
            .O(N__39179),
            .I(measured_delay_hc_23));
    InMux I__8619 (
            .O(N__39174),
            .I(N__39170));
    InMux I__8618 (
            .O(N__39173),
            .I(N__39167));
    LocalMux I__8617 (
            .O(N__39170),
            .I(N__39164));
    LocalMux I__8616 (
            .O(N__39167),
            .I(measured_delay_hc_22));
    Odrv12 I__8615 (
            .O(N__39164),
            .I(measured_delay_hc_22));
    CascadeMux I__8614 (
            .O(N__39159),
            .I(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7Z0Z_19_cascade_ ));
    InMux I__8613 (
            .O(N__39156),
            .I(N__39151));
    InMux I__8612 (
            .O(N__39155),
            .I(N__39148));
    InMux I__8611 (
            .O(N__39154),
            .I(N__39145));
    LocalMux I__8610 (
            .O(N__39151),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__8609 (
            .O(N__39148),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    LocalMux I__8608 (
            .O(N__39145),
            .I(\delay_measurement_inst.delay_hc_reg3lto14 ));
    InMux I__8607 (
            .O(N__39138),
            .I(N__39133));
    InMux I__8606 (
            .O(N__39137),
            .I(N__39130));
    InMux I__8605 (
            .O(N__39136),
            .I(N__39127));
    LocalMux I__8604 (
            .O(N__39133),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__8603 (
            .O(N__39130),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    LocalMux I__8602 (
            .O(N__39127),
            .I(\delay_measurement_inst.delay_hc_reg3lto9 ));
    CascadeMux I__8601 (
            .O(N__39120),
            .I(\delay_measurement_inst.delay_hc_timer.N_299_cascade_ ));
    InMux I__8600 (
            .O(N__39117),
            .I(N__39114));
    LocalMux I__8599 (
            .O(N__39114),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_2_6 ));
    CascadeMux I__8598 (
            .O(N__39111),
            .I(\delay_measurement_inst.N_332_cascade_ ));
    InMux I__8597 (
            .O(N__39108),
            .I(N__39105));
    LocalMux I__8596 (
            .O(N__39105),
            .I(\phase_controller_inst1.stoper_hc.N_406 ));
    CascadeMux I__8595 (
            .O(N__39102),
            .I(\phase_controller_inst1.stoper_hc.N_406_cascade_ ));
    InMux I__8594 (
            .O(N__39099),
            .I(N__39094));
    InMux I__8593 (
            .O(N__39098),
            .I(N__39091));
    InMux I__8592 (
            .O(N__39097),
            .I(N__39088));
    LocalMux I__8591 (
            .O(N__39094),
            .I(N__39085));
    LocalMux I__8590 (
            .O(N__39091),
            .I(N__39082));
    LocalMux I__8589 (
            .O(N__39088),
            .I(N__39079));
    Span4Mux_v I__8588 (
            .O(N__39085),
            .I(N__39075));
    Span4Mux_v I__8587 (
            .O(N__39082),
            .I(N__39070));
    Span4Mux_v I__8586 (
            .O(N__39079),
            .I(N__39070));
    InMux I__8585 (
            .O(N__39078),
            .I(N__39067));
    Odrv4 I__8584 (
            .O(N__39075),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    Odrv4 I__8583 (
            .O(N__39070),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    LocalMux I__8582 (
            .O(N__39067),
            .I(\phase_controller_inst1.stoper_hc.time_passed11 ));
    InMux I__8581 (
            .O(N__39060),
            .I(N__39057));
    LocalMux I__8580 (
            .O(N__39057),
            .I(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_8 ));
    CascadeMux I__8579 (
            .O(N__39054),
            .I(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_7_cascade_ ));
    InMux I__8578 (
            .O(N__39051),
            .I(N__39048));
    LocalMux I__8577 (
            .O(N__39048),
            .I(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_5 ));
    InMux I__8576 (
            .O(N__39045),
            .I(N__39042));
    LocalMux I__8575 (
            .O(N__39042),
            .I(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_6 ));
    CascadeMux I__8574 (
            .O(N__39039),
            .I(N__39036));
    InMux I__8573 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__8572 (
            .O(N__39033),
            .I(N__39030));
    Odrv4 I__8571 (
            .O(N__39030),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__8570 (
            .O(N__39027),
            .I(N__39024));
    InMux I__8569 (
            .O(N__39024),
            .I(N__39021));
    LocalMux I__8568 (
            .O(N__39021),
            .I(N__39018));
    Span4Mux_h I__8567 (
            .O(N__39018),
            .I(N__39015));
    Odrv4 I__8566 (
            .O(N__39015),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__8565 (
            .O(N__39012),
            .I(N__39009));
    InMux I__8564 (
            .O(N__39009),
            .I(N__39006));
    LocalMux I__8563 (
            .O(N__39006),
            .I(N__39003));
    Span4Mux_h I__8562 (
            .O(N__39003),
            .I(N__39000));
    Span4Mux_h I__8561 (
            .O(N__39000),
            .I(N__38997));
    Odrv4 I__8560 (
            .O(N__38997),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__8559 (
            .O(N__38994),
            .I(N__38991));
    InMux I__8558 (
            .O(N__38991),
            .I(N__38988));
    LocalMux I__8557 (
            .O(N__38988),
            .I(N__38985));
    Span4Mux_h I__8556 (
            .O(N__38985),
            .I(N__38982));
    Odrv4 I__8555 (
            .O(N__38982),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__8554 (
            .O(N__38979),
            .I(N__38976));
    InMux I__8553 (
            .O(N__38976),
            .I(N__38973));
    LocalMux I__8552 (
            .O(N__38973),
            .I(N__38970));
    Odrv12 I__8551 (
            .O(N__38970),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__8550 (
            .O(N__38967),
            .I(N__38964));
    InMux I__8549 (
            .O(N__38964),
            .I(N__38961));
    LocalMux I__8548 (
            .O(N__38961),
            .I(N__38958));
    Span4Mux_h I__8547 (
            .O(N__38958),
            .I(N__38955));
    Odrv4 I__8546 (
            .O(N__38955),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__8545 (
            .O(N__38952),
            .I(N__38949));
    InMux I__8544 (
            .O(N__38949),
            .I(N__38946));
    LocalMux I__8543 (
            .O(N__38946),
            .I(N__38943));
    Span4Mux_h I__8542 (
            .O(N__38943),
            .I(N__38940));
    Odrv4 I__8541 (
            .O(N__38940),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CEMux I__8540 (
            .O(N__38937),
            .I(N__38934));
    LocalMux I__8539 (
            .O(N__38934),
            .I(N__38929));
    CEMux I__8538 (
            .O(N__38933),
            .I(N__38926));
    CEMux I__8537 (
            .O(N__38932),
            .I(N__38922));
    Span4Mux_h I__8536 (
            .O(N__38929),
            .I(N__38917));
    LocalMux I__8535 (
            .O(N__38926),
            .I(N__38917));
    CEMux I__8534 (
            .O(N__38925),
            .I(N__38914));
    LocalMux I__8533 (
            .O(N__38922),
            .I(N__38911));
    Span4Mux_v I__8532 (
            .O(N__38917),
            .I(N__38906));
    LocalMux I__8531 (
            .O(N__38914),
            .I(N__38906));
    Span4Mux_v I__8530 (
            .O(N__38911),
            .I(N__38903));
    Span4Mux_h I__8529 (
            .O(N__38906),
            .I(N__38900));
    Span4Mux_v I__8528 (
            .O(N__38903),
            .I(N__38897));
    Span4Mux_v I__8527 (
            .O(N__38900),
            .I(N__38894));
    Odrv4 I__8526 (
            .O(N__38897),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    Odrv4 I__8525 (
            .O(N__38894),
            .I(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ));
    CascadeMux I__8524 (
            .O(N__38889),
            .I(\phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0Z0Z_3_cascade_ ));
    CascadeMux I__8523 (
            .O(N__38886),
            .I(\phase_controller_inst1.stoper_hc.N_316_cascade_ ));
    CascadeMux I__8522 (
            .O(N__38883),
            .I(N__38880));
    InMux I__8521 (
            .O(N__38880),
            .I(N__38877));
    LocalMux I__8520 (
            .O(N__38877),
            .I(N__38874));
    Odrv4 I__8519 (
            .O(N__38874),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ));
    InMux I__8518 (
            .O(N__38871),
            .I(N__38867));
    InMux I__8517 (
            .O(N__38870),
            .I(N__38864));
    LocalMux I__8516 (
            .O(N__38867),
            .I(N__38861));
    LocalMux I__8515 (
            .O(N__38864),
            .I(N__38856));
    Span4Mux_h I__8514 (
            .O(N__38861),
            .I(N__38856));
    Odrv4 I__8513 (
            .O(N__38856),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__8512 (
            .O(N__38853),
            .I(N__38850));
    LocalMux I__8511 (
            .O(N__38850),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ));
    InMux I__8510 (
            .O(N__38847),
            .I(N__38844));
    LocalMux I__8509 (
            .O(N__38844),
            .I(N__38840));
    InMux I__8508 (
            .O(N__38843),
            .I(N__38837));
    Span4Mux_h I__8507 (
            .O(N__38840),
            .I(N__38834));
    LocalMux I__8506 (
            .O(N__38837),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__8505 (
            .O(N__38834),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__8504 (
            .O(N__38829),
            .I(\phase_controller_inst1.stoper_hc.un2_startlt31_5_cascade_ ));
    InMux I__8503 (
            .O(N__38826),
            .I(N__38823));
    LocalMux I__8502 (
            .O(N__38823),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__8501 (
            .O(N__38820),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__8500 (
            .O(N__38817),
            .I(N__38814));
    LocalMux I__8499 (
            .O(N__38814),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__8498 (
            .O(N__38811),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8497 (
            .O(N__38808),
            .I(N__38805));
    InMux I__8496 (
            .O(N__38805),
            .I(N__38802));
    LocalMux I__8495 (
            .O(N__38802),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__8494 (
            .O(N__38799),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__8493 (
            .O(N__38796),
            .I(N__38793));
    LocalMux I__8492 (
            .O(N__38793),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__8491 (
            .O(N__38790),
            .I(bfn_16_14_0_));
    InMux I__8490 (
            .O(N__38787),
            .I(N__38784));
    LocalMux I__8489 (
            .O(N__38784),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__8488 (
            .O(N__38781),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8487 (
            .O(N__38778),
            .I(N__38775));
    LocalMux I__8486 (
            .O(N__38775),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__8485 (
            .O(N__38772),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__8484 (
            .O(N__38769),
            .I(N__38766));
    InMux I__8483 (
            .O(N__38766),
            .I(N__38763));
    LocalMux I__8482 (
            .O(N__38763),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ));
    InMux I__8481 (
            .O(N__38760),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8480 (
            .O(N__38757),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8479 (
            .O(N__38754),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__8478 (
            .O(N__38751),
            .I(N__38746));
    InMux I__8477 (
            .O(N__38750),
            .I(N__38743));
    InMux I__8476 (
            .O(N__38749),
            .I(N__38740));
    LocalMux I__8475 (
            .O(N__38746),
            .I(N__38733));
    LocalMux I__8474 (
            .O(N__38743),
            .I(N__38733));
    LocalMux I__8473 (
            .O(N__38740),
            .I(N__38733));
    Odrv4 I__8472 (
            .O(N__38733),
            .I(\delay_measurement_inst.elapsed_time_tr_16 ));
    InMux I__8471 (
            .O(N__38730),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__8470 (
            .O(N__38727),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__8469 (
            .O(N__38724),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__8468 (
            .O(N__38721),
            .I(N__38716));
    InMux I__8467 (
            .O(N__38720),
            .I(N__38713));
    InMux I__8466 (
            .O(N__38719),
            .I(N__38708));
    InMux I__8465 (
            .O(N__38716),
            .I(N__38708));
    LocalMux I__8464 (
            .O(N__38713),
            .I(N__38705));
    LocalMux I__8463 (
            .O(N__38708),
            .I(N__38702));
    Odrv12 I__8462 (
            .O(N__38705),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    Odrv12 I__8461 (
            .O(N__38702),
            .I(\delay_measurement_inst.elapsed_time_tr_19 ));
    InMux I__8460 (
            .O(N__38697),
            .I(bfn_16_13_0_));
    InMux I__8459 (
            .O(N__38694),
            .I(N__38691));
    LocalMux I__8458 (
            .O(N__38691),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__8457 (
            .O(N__38688),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__8456 (
            .O(N__38685),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8455 (
            .O(N__38682),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__8454 (
            .O(N__38679),
            .I(N__38676));
    LocalMux I__8453 (
            .O(N__38676),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__8452 (
            .O(N__38673),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8451 (
            .O(N__38670),
            .I(N__38667));
    LocalMux I__8450 (
            .O(N__38667),
            .I(N__38664));
    Span4Mux_h I__8449 (
            .O(N__38664),
            .I(N__38660));
    InMux I__8448 (
            .O(N__38663),
            .I(N__38657));
    Odrv4 I__8447 (
            .O(N__38660),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    LocalMux I__8446 (
            .O(N__38657),
            .I(\delay_measurement_inst.elapsed_time_tr_7 ));
    InMux I__8445 (
            .O(N__38652),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__8444 (
            .O(N__38649),
            .I(N__38646));
    LocalMux I__8443 (
            .O(N__38646),
            .I(N__38643));
    Span4Mux_h I__8442 (
            .O(N__38643),
            .I(N__38639));
    InMux I__8441 (
            .O(N__38642),
            .I(N__38636));
    Odrv4 I__8440 (
            .O(N__38639),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    LocalMux I__8439 (
            .O(N__38636),
            .I(\delay_measurement_inst.elapsed_time_tr_8 ));
    InMux I__8438 (
            .O(N__38631),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__8437 (
            .O(N__38628),
            .I(N__38624));
    InMux I__8436 (
            .O(N__38627),
            .I(N__38621));
    LocalMux I__8435 (
            .O(N__38624),
            .I(N__38616));
    LocalMux I__8434 (
            .O(N__38621),
            .I(N__38616));
    Span4Mux_h I__8433 (
            .O(N__38616),
            .I(N__38610));
    InMux I__8432 (
            .O(N__38615),
            .I(N__38607));
    InMux I__8431 (
            .O(N__38614),
            .I(N__38604));
    InMux I__8430 (
            .O(N__38613),
            .I(N__38601));
    Odrv4 I__8429 (
            .O(N__38610),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    LocalMux I__8428 (
            .O(N__38607),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    LocalMux I__8427 (
            .O(N__38604),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    LocalMux I__8426 (
            .O(N__38601),
            .I(\delay_measurement_inst.delay_tr_reg3lto9 ));
    InMux I__8425 (
            .O(N__38592),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__8424 (
            .O(N__38589),
            .I(N__38586));
    LocalMux I__8423 (
            .O(N__38586),
            .I(N__38583));
    Span4Mux_v I__8422 (
            .O(N__38583),
            .I(N__38579));
    InMux I__8421 (
            .O(N__38582),
            .I(N__38576));
    Odrv4 I__8420 (
            .O(N__38579),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    LocalMux I__8419 (
            .O(N__38576),
            .I(\delay_measurement_inst.elapsed_time_tr_10 ));
    InMux I__8418 (
            .O(N__38571),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__8417 (
            .O(N__38568),
            .I(N__38565));
    LocalMux I__8416 (
            .O(N__38565),
            .I(N__38561));
    InMux I__8415 (
            .O(N__38564),
            .I(N__38558));
    Odrv4 I__8414 (
            .O(N__38561),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    LocalMux I__8413 (
            .O(N__38558),
            .I(\delay_measurement_inst.elapsed_time_tr_11 ));
    InMux I__8412 (
            .O(N__38553),
            .I(bfn_16_12_0_));
    InMux I__8411 (
            .O(N__38550),
            .I(N__38547));
    LocalMux I__8410 (
            .O(N__38547),
            .I(N__38543));
    InMux I__8409 (
            .O(N__38546),
            .I(N__38540));
    Odrv4 I__8408 (
            .O(N__38543),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    LocalMux I__8407 (
            .O(N__38540),
            .I(\delay_measurement_inst.elapsed_time_tr_12 ));
    InMux I__8406 (
            .O(N__38535),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__8405 (
            .O(N__38532),
            .I(N__38528));
    CascadeMux I__8404 (
            .O(N__38531),
            .I(N__38525));
    LocalMux I__8403 (
            .O(N__38528),
            .I(N__38522));
    InMux I__8402 (
            .O(N__38525),
            .I(N__38519));
    Odrv4 I__8401 (
            .O(N__38522),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    LocalMux I__8400 (
            .O(N__38519),
            .I(\delay_measurement_inst.elapsed_time_tr_13 ));
    InMux I__8399 (
            .O(N__38514),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__8398 (
            .O(N__38511),
            .I(N__38505));
    InMux I__8397 (
            .O(N__38510),
            .I(N__38502));
    InMux I__8396 (
            .O(N__38509),
            .I(N__38498));
    InMux I__8395 (
            .O(N__38508),
            .I(N__38495));
    LocalMux I__8394 (
            .O(N__38505),
            .I(N__38490));
    LocalMux I__8393 (
            .O(N__38502),
            .I(N__38490));
    InMux I__8392 (
            .O(N__38501),
            .I(N__38487));
    LocalMux I__8391 (
            .O(N__38498),
            .I(N__38484));
    LocalMux I__8390 (
            .O(N__38495),
            .I(N__38481));
    Odrv4 I__8389 (
            .O(N__38490),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    LocalMux I__8388 (
            .O(N__38487),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    Odrv12 I__8387 (
            .O(N__38484),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    Odrv4 I__8386 (
            .O(N__38481),
            .I(\delay_measurement_inst.delay_tr_reg3lto14 ));
    InMux I__8385 (
            .O(N__38472),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__8384 (
            .O(N__38469),
            .I(N__38465));
    CascadeMux I__8383 (
            .O(N__38468),
            .I(N__38461));
    InMux I__8382 (
            .O(N__38465),
            .I(N__38453));
    InMux I__8381 (
            .O(N__38464),
            .I(N__38453));
    InMux I__8380 (
            .O(N__38461),
            .I(N__38448));
    InMux I__8379 (
            .O(N__38460),
            .I(N__38443));
    InMux I__8378 (
            .O(N__38459),
            .I(N__38443));
    CascadeMux I__8377 (
            .O(N__38458),
            .I(N__38439));
    LocalMux I__8376 (
            .O(N__38453),
            .I(N__38436));
    InMux I__8375 (
            .O(N__38452),
            .I(N__38431));
    InMux I__8374 (
            .O(N__38451),
            .I(N__38431));
    LocalMux I__8373 (
            .O(N__38448),
            .I(N__38428));
    LocalMux I__8372 (
            .O(N__38443),
            .I(N__38425));
    InMux I__8371 (
            .O(N__38442),
            .I(N__38420));
    InMux I__8370 (
            .O(N__38439),
            .I(N__38420));
    Span4Mux_v I__8369 (
            .O(N__38436),
            .I(N__38415));
    LocalMux I__8368 (
            .O(N__38431),
            .I(N__38415));
    Span4Mux_h I__8367 (
            .O(N__38428),
            .I(N__38412));
    Odrv4 I__8366 (
            .O(N__38425),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    LocalMux I__8365 (
            .O(N__38420),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv4 I__8364 (
            .O(N__38415),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    Odrv4 I__8363 (
            .O(N__38412),
            .I(\delay_measurement_inst.delay_tr_reg3lto15 ));
    InMux I__8362 (
            .O(N__38403),
            .I(N__38398));
    InMux I__8361 (
            .O(N__38402),
            .I(N__38395));
    InMux I__8360 (
            .O(N__38401),
            .I(N__38392));
    LocalMux I__8359 (
            .O(N__38398),
            .I(N__38389));
    LocalMux I__8358 (
            .O(N__38395),
            .I(N__38386));
    LocalMux I__8357 (
            .O(N__38392),
            .I(N__38381));
    Span4Mux_v I__8356 (
            .O(N__38389),
            .I(N__38381));
    Odrv12 I__8355 (
            .O(N__38386),
            .I(il_min_comp1_D2));
    Odrv4 I__8354 (
            .O(N__38381),
            .I(il_min_comp1_D2));
    InMux I__8353 (
            .O(N__38376),
            .I(N__38373));
    LocalMux I__8352 (
            .O(N__38373),
            .I(N__38370));
    Odrv4 I__8351 (
            .O(N__38370),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__8350 (
            .O(N__38367),
            .I(N__38364));
    LocalMux I__8349 (
            .O(N__38364),
            .I(N__38360));
    InMux I__8348 (
            .O(N__38363),
            .I(N__38357));
    Span4Mux_v I__8347 (
            .O(N__38360),
            .I(N__38351));
    LocalMux I__8346 (
            .O(N__38357),
            .I(N__38351));
    InMux I__8345 (
            .O(N__38356),
            .I(N__38348));
    Span4Mux_v I__8344 (
            .O(N__38351),
            .I(N__38345));
    LocalMux I__8343 (
            .O(N__38348),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    Odrv4 I__8342 (
            .O(N__38345),
            .I(\delay_measurement_inst.elapsed_time_tr_2 ));
    CascadeMux I__8341 (
            .O(N__38340),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ));
    InMux I__8340 (
            .O(N__38337),
            .I(N__38334));
    LocalMux I__8339 (
            .O(N__38334),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ));
    InMux I__8338 (
            .O(N__38331),
            .I(N__38325));
    InMux I__8337 (
            .O(N__38330),
            .I(N__38325));
    LocalMux I__8336 (
            .O(N__38325),
            .I(\delay_measurement_inst.delay_tr_timer.N_373_4 ));
    InMux I__8335 (
            .O(N__38322),
            .I(N__38319));
    LocalMux I__8334 (
            .O(N__38319),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ));
    InMux I__8333 (
            .O(N__38316),
            .I(N__38313));
    LocalMux I__8332 (
            .O(N__38313),
            .I(N__38308));
    InMux I__8331 (
            .O(N__38312),
            .I(N__38303));
    InMux I__8330 (
            .O(N__38311),
            .I(N__38303));
    Odrv4 I__8329 (
            .O(N__38308),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    LocalMux I__8328 (
            .O(N__38303),
            .I(\delay_measurement_inst.elapsed_time_tr_3 ));
    InMux I__8327 (
            .O(N__38298),
            .I(N__38295));
    LocalMux I__8326 (
            .O(N__38295),
            .I(N__38291));
    InMux I__8325 (
            .O(N__38294),
            .I(N__38288));
    Odrv4 I__8324 (
            .O(N__38291),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    LocalMux I__8323 (
            .O(N__38288),
            .I(\delay_measurement_inst.elapsed_time_tr_4 ));
    InMux I__8322 (
            .O(N__38283),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__8321 (
            .O(N__38280),
            .I(N__38277));
    LocalMux I__8320 (
            .O(N__38277),
            .I(N__38273));
    InMux I__8319 (
            .O(N__38276),
            .I(N__38270));
    Odrv4 I__8318 (
            .O(N__38273),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    LocalMux I__8317 (
            .O(N__38270),
            .I(\delay_measurement_inst.elapsed_time_tr_5 ));
    InMux I__8316 (
            .O(N__38265),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__8315 (
            .O(N__38262),
            .I(N__38256));
    InMux I__8314 (
            .O(N__38261),
            .I(N__38253));
    InMux I__8313 (
            .O(N__38260),
            .I(N__38250));
    InMux I__8312 (
            .O(N__38259),
            .I(N__38247));
    LocalMux I__8311 (
            .O(N__38256),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    LocalMux I__8310 (
            .O(N__38253),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    LocalMux I__8309 (
            .O(N__38250),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    LocalMux I__8308 (
            .O(N__38247),
            .I(\delay_measurement_inst.delay_tr_reg3lto6 ));
    InMux I__8307 (
            .O(N__38238),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__8306 (
            .O(N__38235),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_ ));
    InMux I__8305 (
            .O(N__38232),
            .I(N__38227));
    InMux I__8304 (
            .O(N__38231),
            .I(N__38224));
    InMux I__8303 (
            .O(N__38230),
            .I(N__38221));
    LocalMux I__8302 (
            .O(N__38227),
            .I(N__38218));
    LocalMux I__8301 (
            .O(N__38224),
            .I(N__38214));
    LocalMux I__8300 (
            .O(N__38221),
            .I(N__38210));
    Span4Mux_v I__8299 (
            .O(N__38218),
            .I(N__38207));
    InMux I__8298 (
            .O(N__38217),
            .I(N__38204));
    Span4Mux_h I__8297 (
            .O(N__38214),
            .I(N__38201));
    InMux I__8296 (
            .O(N__38213),
            .I(N__38198));
    Span4Mux_v I__8295 (
            .O(N__38210),
            .I(N__38195));
    Span4Mux_h I__8294 (
            .O(N__38207),
            .I(N__38190));
    LocalMux I__8293 (
            .O(N__38204),
            .I(N__38190));
    Span4Mux_h I__8292 (
            .O(N__38201),
            .I(N__38187));
    LocalMux I__8291 (
            .O(N__38198),
            .I(N__38183));
    Span4Mux_h I__8290 (
            .O(N__38195),
            .I(N__38178));
    Span4Mux_v I__8289 (
            .O(N__38190),
            .I(N__38178));
    Sp12to4 I__8288 (
            .O(N__38187),
            .I(N__38175));
    InMux I__8287 (
            .O(N__38186),
            .I(N__38172));
    Span4Mux_v I__8286 (
            .O(N__38183),
            .I(N__38167));
    Span4Mux_h I__8285 (
            .O(N__38178),
            .I(N__38167));
    Odrv12 I__8284 (
            .O(N__38175),
            .I(phase_controller_inst1_state_4));
    LocalMux I__8283 (
            .O(N__38172),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__8282 (
            .O(N__38167),
            .I(phase_controller_inst1_state_4));
    InMux I__8281 (
            .O(N__38160),
            .I(N__38157));
    LocalMux I__8280 (
            .O(N__38157),
            .I(N__38153));
    InMux I__8279 (
            .O(N__38156),
            .I(N__38150));
    Span4Mux_h I__8278 (
            .O(N__38153),
            .I(N__38146));
    LocalMux I__8277 (
            .O(N__38150),
            .I(N__38143));
    InMux I__8276 (
            .O(N__38149),
            .I(N__38140));
    Odrv4 I__8275 (
            .O(N__38146),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    Odrv12 I__8274 (
            .O(N__38143),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    LocalMux I__8273 (
            .O(N__38140),
            .I(\phase_controller_inst1.stoper_tr.time_passed11 ));
    CascadeMux I__8272 (
            .O(N__38133),
            .I(N__38130));
    InMux I__8271 (
            .O(N__38130),
            .I(N__38127));
    LocalMux I__8270 (
            .O(N__38127),
            .I(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ));
    InMux I__8269 (
            .O(N__38124),
            .I(N__38121));
    LocalMux I__8268 (
            .O(N__38121),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ));
    InMux I__8267 (
            .O(N__38118),
            .I(N__38115));
    LocalMux I__8266 (
            .O(N__38115),
            .I(N__38111));
    InMux I__8265 (
            .O(N__38114),
            .I(N__38108));
    Span4Mux_v I__8264 (
            .O(N__38111),
            .I(N__38105));
    LocalMux I__8263 (
            .O(N__38108),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8262 (
            .O(N__38105),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__8261 (
            .O(N__38100),
            .I(N__38096));
    InMux I__8260 (
            .O(N__38099),
            .I(N__38088));
    InMux I__8259 (
            .O(N__38096),
            .I(N__38088));
    InMux I__8258 (
            .O(N__38095),
            .I(N__38088));
    LocalMux I__8257 (
            .O(N__38088),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__8256 (
            .O(N__38085),
            .I(N__38079));
    InMux I__8255 (
            .O(N__38084),
            .I(N__38079));
    LocalMux I__8254 (
            .O(N__38079),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__8253 (
            .O(N__38076),
            .I(N__38070));
    InMux I__8252 (
            .O(N__38075),
            .I(N__38067));
    InMux I__8251 (
            .O(N__38074),
            .I(N__38062));
    InMux I__8250 (
            .O(N__38073),
            .I(N__38062));
    LocalMux I__8249 (
            .O(N__38070),
            .I(N__38059));
    LocalMux I__8248 (
            .O(N__38067),
            .I(N__38054));
    LocalMux I__8247 (
            .O(N__38062),
            .I(N__38054));
    Span12Mux_h I__8246 (
            .O(N__38059),
            .I(N__38051));
    Span4Mux_h I__8245 (
            .O(N__38054),
            .I(N__38048));
    Odrv12 I__8244 (
            .O(N__38051),
            .I(measured_delay_tr_16));
    Odrv4 I__8243 (
            .O(N__38048),
            .I(measured_delay_tr_16));
    InMux I__8242 (
            .O(N__38043),
            .I(N__38038));
    CascadeMux I__8241 (
            .O(N__38042),
            .I(N__38034));
    CascadeMux I__8240 (
            .O(N__38041),
            .I(N__38031));
    LocalMux I__8239 (
            .O(N__38038),
            .I(N__38028));
    InMux I__8238 (
            .O(N__38037),
            .I(N__38025));
    InMux I__8237 (
            .O(N__38034),
            .I(N__38020));
    InMux I__8236 (
            .O(N__38031),
            .I(N__38020));
    Span4Mux_v I__8235 (
            .O(N__38028),
            .I(N__38017));
    LocalMux I__8234 (
            .O(N__38025),
            .I(N__38014));
    LocalMux I__8233 (
            .O(N__38020),
            .I(N__38011));
    Span4Mux_h I__8232 (
            .O(N__38017),
            .I(N__38008));
    Span4Mux_h I__8231 (
            .O(N__38014),
            .I(N__38005));
    Span4Mux_h I__8230 (
            .O(N__38011),
            .I(N__38002));
    Odrv4 I__8229 (
            .O(N__38008),
            .I(measured_delay_tr_19));
    Odrv4 I__8228 (
            .O(N__38005),
            .I(measured_delay_tr_19));
    Odrv4 I__8227 (
            .O(N__38002),
            .I(measured_delay_tr_19));
    CascadeMux I__8226 (
            .O(N__37995),
            .I(N__37990));
    InMux I__8225 (
            .O(N__37994),
            .I(N__37985));
    InMux I__8224 (
            .O(N__37993),
            .I(N__37985));
    InMux I__8223 (
            .O(N__37990),
            .I(N__37982));
    LocalMux I__8222 (
            .O(N__37985),
            .I(N__37977));
    LocalMux I__8221 (
            .O(N__37982),
            .I(N__37977));
    Span4Mux_h I__8220 (
            .O(N__37977),
            .I(N__37973));
    InMux I__8219 (
            .O(N__37976),
            .I(N__37970));
    Odrv4 I__8218 (
            .O(N__37973),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ));
    LocalMux I__8217 (
            .O(N__37970),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ));
    CascadeMux I__8216 (
            .O(N__37965),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16_cascade_ ));
    InMux I__8215 (
            .O(N__37962),
            .I(N__37959));
    LocalMux I__8214 (
            .O(N__37959),
            .I(N__37956));
    Odrv12 I__8213 (
            .O(N__37956),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_2 ));
    InMux I__8212 (
            .O(N__37953),
            .I(N__37950));
    LocalMux I__8211 (
            .O(N__37950),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_6 ));
    InMux I__8210 (
            .O(N__37947),
            .I(N__37942));
    InMux I__8209 (
            .O(N__37946),
            .I(N__37939));
    InMux I__8208 (
            .O(N__37945),
            .I(N__37936));
    LocalMux I__8207 (
            .O(N__37942),
            .I(N__37933));
    LocalMux I__8206 (
            .O(N__37939),
            .I(N__37929));
    LocalMux I__8205 (
            .O(N__37936),
            .I(N__37926));
    Span4Mux_v I__8204 (
            .O(N__37933),
            .I(N__37923));
    InMux I__8203 (
            .O(N__37932),
            .I(N__37920));
    Span4Mux_h I__8202 (
            .O(N__37929),
            .I(N__37917));
    Odrv4 I__8201 (
            .O(N__37926),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__8200 (
            .O(N__37923),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__8199 (
            .O(N__37920),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__8198 (
            .O(N__37917),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    InMux I__8197 (
            .O(N__37908),
            .I(N__37905));
    LocalMux I__8196 (
            .O(N__37905),
            .I(N__37901));
    InMux I__8195 (
            .O(N__37904),
            .I(N__37898));
    Span4Mux_v I__8194 (
            .O(N__37901),
            .I(N__37895));
    LocalMux I__8193 (
            .O(N__37898),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__8192 (
            .O(N__37895),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__8191 (
            .O(N__37890),
            .I(N__37886));
    CascadeMux I__8190 (
            .O(N__37889),
            .I(N__37883));
    InMux I__8189 (
            .O(N__37886),
            .I(N__37877));
    InMux I__8188 (
            .O(N__37883),
            .I(N__37877));
    InMux I__8187 (
            .O(N__37882),
            .I(N__37874));
    LocalMux I__8186 (
            .O(N__37877),
            .I(N__37871));
    LocalMux I__8185 (
            .O(N__37874),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__8184 (
            .O(N__37871),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__8183 (
            .O(N__37866),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8182 (
            .O(N__37863),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__8181 (
            .O(N__37860),
            .I(N__37845));
    CEMux I__8180 (
            .O(N__37859),
            .I(N__37845));
    CEMux I__8179 (
            .O(N__37858),
            .I(N__37845));
    CEMux I__8178 (
            .O(N__37857),
            .I(N__37845));
    CEMux I__8177 (
            .O(N__37856),
            .I(N__37845));
    GlobalMux I__8176 (
            .O(N__37845),
            .I(N__37842));
    gio2CtrlBuf I__8175 (
            .O(N__37842),
            .I(\delay_measurement_inst.delay_hc_timer.N_461_i_g ));
    InMux I__8174 (
            .O(N__37839),
            .I(N__37835));
    InMux I__8173 (
            .O(N__37838),
            .I(N__37832));
    LocalMux I__8172 (
            .O(N__37835),
            .I(N__37829));
    LocalMux I__8171 (
            .O(N__37832),
            .I(N__37826));
    Span12Mux_v I__8170 (
            .O(N__37829),
            .I(N__37823));
    Odrv4 I__8169 (
            .O(N__37826),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv12 I__8168 (
            .O(N__37823),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    CEMux I__8167 (
            .O(N__37818),
            .I(N__37815));
    LocalMux I__8166 (
            .O(N__37815),
            .I(N__37812));
    Span4Mux_v I__8165 (
            .O(N__37812),
            .I(N__37806));
    CEMux I__8164 (
            .O(N__37811),
            .I(N__37803));
    CEMux I__8163 (
            .O(N__37810),
            .I(N__37800));
    CEMux I__8162 (
            .O(N__37809),
            .I(N__37797));
    Span4Mux_h I__8161 (
            .O(N__37806),
            .I(N__37792));
    LocalMux I__8160 (
            .O(N__37803),
            .I(N__37792));
    LocalMux I__8159 (
            .O(N__37800),
            .I(N__37787));
    LocalMux I__8158 (
            .O(N__37797),
            .I(N__37787));
    Span4Mux_h I__8157 (
            .O(N__37792),
            .I(N__37784));
    Odrv4 I__8156 (
            .O(N__37787),
            .I(\delay_measurement_inst.delay_hc_timer.N_462_i ));
    Odrv4 I__8155 (
            .O(N__37784),
            .I(\delay_measurement_inst.delay_hc_timer.N_462_i ));
    InMux I__8154 (
            .O(N__37779),
            .I(N__37755));
    InMux I__8153 (
            .O(N__37778),
            .I(N__37755));
    InMux I__8152 (
            .O(N__37777),
            .I(N__37755));
    InMux I__8151 (
            .O(N__37776),
            .I(N__37755));
    InMux I__8150 (
            .O(N__37775),
            .I(N__37746));
    InMux I__8149 (
            .O(N__37774),
            .I(N__37746));
    InMux I__8148 (
            .O(N__37773),
            .I(N__37746));
    InMux I__8147 (
            .O(N__37772),
            .I(N__37746));
    InMux I__8146 (
            .O(N__37771),
            .I(N__37737));
    InMux I__8145 (
            .O(N__37770),
            .I(N__37737));
    InMux I__8144 (
            .O(N__37769),
            .I(N__37737));
    InMux I__8143 (
            .O(N__37768),
            .I(N__37737));
    InMux I__8142 (
            .O(N__37767),
            .I(N__37714));
    InMux I__8141 (
            .O(N__37766),
            .I(N__37714));
    InMux I__8140 (
            .O(N__37765),
            .I(N__37714));
    InMux I__8139 (
            .O(N__37764),
            .I(N__37714));
    LocalMux I__8138 (
            .O(N__37755),
            .I(N__37709));
    LocalMux I__8137 (
            .O(N__37746),
            .I(N__37709));
    LocalMux I__8136 (
            .O(N__37737),
            .I(N__37706));
    InMux I__8135 (
            .O(N__37736),
            .I(N__37697));
    InMux I__8134 (
            .O(N__37735),
            .I(N__37697));
    InMux I__8133 (
            .O(N__37734),
            .I(N__37697));
    InMux I__8132 (
            .O(N__37733),
            .I(N__37697));
    InMux I__8131 (
            .O(N__37732),
            .I(N__37692));
    InMux I__8130 (
            .O(N__37731),
            .I(N__37692));
    InMux I__8129 (
            .O(N__37730),
            .I(N__37683));
    InMux I__8128 (
            .O(N__37729),
            .I(N__37683));
    InMux I__8127 (
            .O(N__37728),
            .I(N__37683));
    InMux I__8126 (
            .O(N__37727),
            .I(N__37683));
    InMux I__8125 (
            .O(N__37726),
            .I(N__37674));
    InMux I__8124 (
            .O(N__37725),
            .I(N__37674));
    InMux I__8123 (
            .O(N__37724),
            .I(N__37674));
    InMux I__8122 (
            .O(N__37723),
            .I(N__37674));
    LocalMux I__8121 (
            .O(N__37714),
            .I(N__37669));
    Span4Mux_v I__8120 (
            .O(N__37709),
            .I(N__37669));
    Span4Mux_h I__8119 (
            .O(N__37706),
            .I(N__37666));
    LocalMux I__8118 (
            .O(N__37697),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__8117 (
            .O(N__37692),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__8116 (
            .O(N__37683),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__8115 (
            .O(N__37674),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8114 (
            .O(N__37669),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8113 (
            .O(N__37666),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__8112 (
            .O(N__37653),
            .I(N__37650));
    LocalMux I__8111 (
            .O(N__37650),
            .I(N__37645));
    InMux I__8110 (
            .O(N__37649),
            .I(N__37641));
    InMux I__8109 (
            .O(N__37648),
            .I(N__37638));
    Span4Mux_v I__8108 (
            .O(N__37645),
            .I(N__37635));
    InMux I__8107 (
            .O(N__37644),
            .I(N__37632));
    LocalMux I__8106 (
            .O(N__37641),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__8105 (
            .O(N__37638),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__8104 (
            .O(N__37635),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__8103 (
            .O(N__37632),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__8102 (
            .O(N__37623),
            .I(N__37620));
    LocalMux I__8101 (
            .O(N__37620),
            .I(N__37617));
    Span12Mux_v I__8100 (
            .O(N__37617),
            .I(N__37614));
    Odrv12 I__8099 (
            .O(N__37614),
            .I(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ));
    InMux I__8098 (
            .O(N__37611),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__8097 (
            .O(N__37608),
            .I(N__37604));
    CascadeMux I__8096 (
            .O(N__37607),
            .I(N__37601));
    InMux I__8095 (
            .O(N__37604),
            .I(N__37596));
    InMux I__8094 (
            .O(N__37601),
            .I(N__37596));
    LocalMux I__8093 (
            .O(N__37596),
            .I(N__37592));
    InMux I__8092 (
            .O(N__37595),
            .I(N__37589));
    Span4Mux_h I__8091 (
            .O(N__37592),
            .I(N__37586));
    LocalMux I__8090 (
            .O(N__37589),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__8089 (
            .O(N__37586),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__8088 (
            .O(N__37581),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__8087 (
            .O(N__37578),
            .I(N__37572));
    InMux I__8086 (
            .O(N__37577),
            .I(N__37572));
    LocalMux I__8085 (
            .O(N__37572),
            .I(N__37568));
    InMux I__8084 (
            .O(N__37571),
            .I(N__37565));
    Span4Mux_v I__8083 (
            .O(N__37568),
            .I(N__37562));
    LocalMux I__8082 (
            .O(N__37565),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__8081 (
            .O(N__37562),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__8080 (
            .O(N__37557),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8079 (
            .O(N__37554),
            .I(N__37548));
    InMux I__8078 (
            .O(N__37553),
            .I(N__37548));
    LocalMux I__8077 (
            .O(N__37548),
            .I(N__37544));
    InMux I__8076 (
            .O(N__37547),
            .I(N__37541));
    Span4Mux_v I__8075 (
            .O(N__37544),
            .I(N__37538));
    LocalMux I__8074 (
            .O(N__37541),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__8073 (
            .O(N__37538),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__8072 (
            .O(N__37533),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__8071 (
            .O(N__37530),
            .I(N__37526));
    CascadeMux I__8070 (
            .O(N__37529),
            .I(N__37523));
    InMux I__8069 (
            .O(N__37526),
            .I(N__37518));
    InMux I__8068 (
            .O(N__37523),
            .I(N__37518));
    LocalMux I__8067 (
            .O(N__37518),
            .I(N__37514));
    InMux I__8066 (
            .O(N__37517),
            .I(N__37511));
    Span4Mux_h I__8065 (
            .O(N__37514),
            .I(N__37508));
    LocalMux I__8064 (
            .O(N__37511),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__8063 (
            .O(N__37508),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__8062 (
            .O(N__37503),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__8061 (
            .O(N__37500),
            .I(N__37496));
    CascadeMux I__8060 (
            .O(N__37499),
            .I(N__37493));
    InMux I__8059 (
            .O(N__37496),
            .I(N__37488));
    InMux I__8058 (
            .O(N__37493),
            .I(N__37488));
    LocalMux I__8057 (
            .O(N__37488),
            .I(N__37484));
    InMux I__8056 (
            .O(N__37487),
            .I(N__37481));
    Span4Mux_h I__8055 (
            .O(N__37484),
            .I(N__37478));
    LocalMux I__8054 (
            .O(N__37481),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__8053 (
            .O(N__37478),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__8052 (
            .O(N__37473),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__8051 (
            .O(N__37470),
            .I(N__37466));
    InMux I__8050 (
            .O(N__37469),
            .I(N__37463));
    LocalMux I__8049 (
            .O(N__37466),
            .I(N__37459));
    LocalMux I__8048 (
            .O(N__37463),
            .I(N__37456));
    InMux I__8047 (
            .O(N__37462),
            .I(N__37453));
    Span4Mux_h I__8046 (
            .O(N__37459),
            .I(N__37450));
    Odrv4 I__8045 (
            .O(N__37456),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__8044 (
            .O(N__37453),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__8043 (
            .O(N__37450),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__8042 (
            .O(N__37443),
            .I(bfn_15_25_0_));
    InMux I__8041 (
            .O(N__37440),
            .I(N__37436));
    InMux I__8040 (
            .O(N__37439),
            .I(N__37433));
    LocalMux I__8039 (
            .O(N__37436),
            .I(N__37429));
    LocalMux I__8038 (
            .O(N__37433),
            .I(N__37426));
    InMux I__8037 (
            .O(N__37432),
            .I(N__37423));
    Span4Mux_h I__8036 (
            .O(N__37429),
            .I(N__37420));
    Odrv4 I__8035 (
            .O(N__37426),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__8034 (
            .O(N__37423),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__8033 (
            .O(N__37420),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__8032 (
            .O(N__37413),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8031 (
            .O(N__37410),
            .I(N__37407));
    LocalMux I__8030 (
            .O(N__37407),
            .I(N__37403));
    InMux I__8029 (
            .O(N__37406),
            .I(N__37400));
    Span4Mux_v I__8028 (
            .O(N__37403),
            .I(N__37397));
    LocalMux I__8027 (
            .O(N__37400),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__8026 (
            .O(N__37397),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__8025 (
            .O(N__37392),
            .I(N__37388));
    CascadeMux I__8024 (
            .O(N__37391),
            .I(N__37385));
    InMux I__8023 (
            .O(N__37388),
            .I(N__37379));
    InMux I__8022 (
            .O(N__37385),
            .I(N__37379));
    InMux I__8021 (
            .O(N__37384),
            .I(N__37376));
    LocalMux I__8020 (
            .O(N__37379),
            .I(N__37373));
    LocalMux I__8019 (
            .O(N__37376),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__8018 (
            .O(N__37373),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__8017 (
            .O(N__37368),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__8016 (
            .O(N__37365),
            .I(N__37361));
    CascadeMux I__8015 (
            .O(N__37364),
            .I(N__37358));
    InMux I__8014 (
            .O(N__37361),
            .I(N__37352));
    InMux I__8013 (
            .O(N__37358),
            .I(N__37352));
    InMux I__8012 (
            .O(N__37357),
            .I(N__37349));
    LocalMux I__8011 (
            .O(N__37352),
            .I(N__37346));
    LocalMux I__8010 (
            .O(N__37349),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__8009 (
            .O(N__37346),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__8008 (
            .O(N__37341),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__8007 (
            .O(N__37338),
            .I(N__37334));
    CascadeMux I__8006 (
            .O(N__37337),
            .I(N__37331));
    InMux I__8005 (
            .O(N__37334),
            .I(N__37326));
    InMux I__8004 (
            .O(N__37331),
            .I(N__37326));
    LocalMux I__8003 (
            .O(N__37326),
            .I(N__37322));
    InMux I__8002 (
            .O(N__37325),
            .I(N__37319));
    Span4Mux_h I__8001 (
            .O(N__37322),
            .I(N__37316));
    LocalMux I__8000 (
            .O(N__37319),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__7999 (
            .O(N__37316),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__7998 (
            .O(N__37311),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__7997 (
            .O(N__37308),
            .I(N__37301));
    InMux I__7996 (
            .O(N__37307),
            .I(N__37301));
    InMux I__7995 (
            .O(N__37306),
            .I(N__37298));
    LocalMux I__7994 (
            .O(N__37301),
            .I(N__37295));
    LocalMux I__7993 (
            .O(N__37298),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__7992 (
            .O(N__37295),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__7991 (
            .O(N__37290),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__7990 (
            .O(N__37287),
            .I(N__37281));
    InMux I__7989 (
            .O(N__37286),
            .I(N__37281));
    LocalMux I__7988 (
            .O(N__37281),
            .I(N__37277));
    InMux I__7987 (
            .O(N__37280),
            .I(N__37274));
    Span4Mux_v I__7986 (
            .O(N__37277),
            .I(N__37271));
    LocalMux I__7985 (
            .O(N__37274),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__7984 (
            .O(N__37271),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__7983 (
            .O(N__37266),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7982 (
            .O(N__37263),
            .I(N__37259));
    CascadeMux I__7981 (
            .O(N__37262),
            .I(N__37256));
    InMux I__7980 (
            .O(N__37259),
            .I(N__37251));
    InMux I__7979 (
            .O(N__37256),
            .I(N__37251));
    LocalMux I__7978 (
            .O(N__37251),
            .I(N__37247));
    InMux I__7977 (
            .O(N__37250),
            .I(N__37244));
    Span4Mux_h I__7976 (
            .O(N__37247),
            .I(N__37241));
    LocalMux I__7975 (
            .O(N__37244),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__7974 (
            .O(N__37241),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__7973 (
            .O(N__37236),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__7972 (
            .O(N__37233),
            .I(N__37229));
    CascadeMux I__7971 (
            .O(N__37232),
            .I(N__37226));
    InMux I__7970 (
            .O(N__37229),
            .I(N__37221));
    InMux I__7969 (
            .O(N__37226),
            .I(N__37221));
    LocalMux I__7968 (
            .O(N__37221),
            .I(N__37217));
    InMux I__7967 (
            .O(N__37220),
            .I(N__37214));
    Span4Mux_h I__7966 (
            .O(N__37217),
            .I(N__37211));
    LocalMux I__7965 (
            .O(N__37214),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__7964 (
            .O(N__37211),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__7963 (
            .O(N__37206),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__7962 (
            .O(N__37203),
            .I(N__37199));
    InMux I__7961 (
            .O(N__37202),
            .I(N__37196));
    LocalMux I__7960 (
            .O(N__37199),
            .I(N__37192));
    LocalMux I__7959 (
            .O(N__37196),
            .I(N__37189));
    InMux I__7958 (
            .O(N__37195),
            .I(N__37186));
    Span4Mux_h I__7957 (
            .O(N__37192),
            .I(N__37183));
    Odrv4 I__7956 (
            .O(N__37189),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__7955 (
            .O(N__37186),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__7954 (
            .O(N__37183),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__7953 (
            .O(N__37176),
            .I(bfn_15_24_0_));
    InMux I__7952 (
            .O(N__37173),
            .I(N__37169));
    InMux I__7951 (
            .O(N__37172),
            .I(N__37166));
    LocalMux I__7950 (
            .O(N__37169),
            .I(N__37162));
    LocalMux I__7949 (
            .O(N__37166),
            .I(N__37159));
    InMux I__7948 (
            .O(N__37165),
            .I(N__37156));
    Span4Mux_h I__7947 (
            .O(N__37162),
            .I(N__37153));
    Odrv4 I__7946 (
            .O(N__37159),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__7945 (
            .O(N__37156),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__7944 (
            .O(N__37153),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__7943 (
            .O(N__37146),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__7942 (
            .O(N__37143),
            .I(N__37139));
    CascadeMux I__7941 (
            .O(N__37142),
            .I(N__37136));
    InMux I__7940 (
            .O(N__37139),
            .I(N__37130));
    InMux I__7939 (
            .O(N__37136),
            .I(N__37130));
    InMux I__7938 (
            .O(N__37135),
            .I(N__37127));
    LocalMux I__7937 (
            .O(N__37130),
            .I(N__37124));
    LocalMux I__7936 (
            .O(N__37127),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__7935 (
            .O(N__37124),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    CascadeMux I__7934 (
            .O(N__37119),
            .I(N__37115));
    CascadeMux I__7933 (
            .O(N__37118),
            .I(N__37112));
    InMux I__7932 (
            .O(N__37115),
            .I(N__37106));
    InMux I__7931 (
            .O(N__37112),
            .I(N__37106));
    InMux I__7930 (
            .O(N__37111),
            .I(N__37103));
    LocalMux I__7929 (
            .O(N__37106),
            .I(N__37100));
    LocalMux I__7928 (
            .O(N__37103),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__7927 (
            .O(N__37100),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__7926 (
            .O(N__37095),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__7925 (
            .O(N__37092),
            .I(N__37088));
    CascadeMux I__7924 (
            .O(N__37091),
            .I(N__37085));
    InMux I__7923 (
            .O(N__37088),
            .I(N__37080));
    InMux I__7922 (
            .O(N__37085),
            .I(N__37080));
    LocalMux I__7921 (
            .O(N__37080),
            .I(N__37076));
    InMux I__7920 (
            .O(N__37079),
            .I(N__37073));
    Span4Mux_h I__7919 (
            .O(N__37076),
            .I(N__37070));
    LocalMux I__7918 (
            .O(N__37073),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__7917 (
            .O(N__37070),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__7916 (
            .O(N__37065),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__7915 (
            .O(N__37062),
            .I(N__37056));
    InMux I__7914 (
            .O(N__37061),
            .I(N__37056));
    LocalMux I__7913 (
            .O(N__37056),
            .I(N__37052));
    InMux I__7912 (
            .O(N__37055),
            .I(N__37049));
    Span4Mux_v I__7911 (
            .O(N__37052),
            .I(N__37046));
    LocalMux I__7910 (
            .O(N__37049),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__7909 (
            .O(N__37046),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__7908 (
            .O(N__37041),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__7907 (
            .O(N__37038),
            .I(N__37032));
    InMux I__7906 (
            .O(N__37037),
            .I(N__37032));
    LocalMux I__7905 (
            .O(N__37032),
            .I(N__37028));
    InMux I__7904 (
            .O(N__37031),
            .I(N__37025));
    Span4Mux_v I__7903 (
            .O(N__37028),
            .I(N__37022));
    LocalMux I__7902 (
            .O(N__37025),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__7901 (
            .O(N__37022),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__7900 (
            .O(N__37017),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7899 (
            .O(N__37014),
            .I(N__37010));
    CascadeMux I__7898 (
            .O(N__37013),
            .I(N__37007));
    InMux I__7897 (
            .O(N__37010),
            .I(N__37002));
    InMux I__7896 (
            .O(N__37007),
            .I(N__37002));
    LocalMux I__7895 (
            .O(N__37002),
            .I(N__36998));
    InMux I__7894 (
            .O(N__37001),
            .I(N__36995));
    Span4Mux_h I__7893 (
            .O(N__36998),
            .I(N__36992));
    LocalMux I__7892 (
            .O(N__36995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__7891 (
            .O(N__36992),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__7890 (
            .O(N__36987),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__7889 (
            .O(N__36984),
            .I(N__36980));
    CascadeMux I__7888 (
            .O(N__36983),
            .I(N__36977));
    InMux I__7887 (
            .O(N__36980),
            .I(N__36972));
    InMux I__7886 (
            .O(N__36977),
            .I(N__36972));
    LocalMux I__7885 (
            .O(N__36972),
            .I(N__36968));
    InMux I__7884 (
            .O(N__36971),
            .I(N__36965));
    Span4Mux_h I__7883 (
            .O(N__36968),
            .I(N__36962));
    LocalMux I__7882 (
            .O(N__36965),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__7881 (
            .O(N__36962),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__7880 (
            .O(N__36957),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__7879 (
            .O(N__36954),
            .I(N__36950));
    InMux I__7878 (
            .O(N__36953),
            .I(N__36947));
    LocalMux I__7877 (
            .O(N__36950),
            .I(N__36944));
    LocalMux I__7876 (
            .O(N__36947),
            .I(N__36940));
    Span4Mux_h I__7875 (
            .O(N__36944),
            .I(N__36937));
    InMux I__7874 (
            .O(N__36943),
            .I(N__36934));
    Span4Mux_h I__7873 (
            .O(N__36940),
            .I(N__36931));
    Odrv4 I__7872 (
            .O(N__36937),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__7871 (
            .O(N__36934),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__7870 (
            .O(N__36931),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__7869 (
            .O(N__36924),
            .I(bfn_15_23_0_));
    InMux I__7868 (
            .O(N__36921),
            .I(N__36917));
    InMux I__7867 (
            .O(N__36920),
            .I(N__36914));
    LocalMux I__7866 (
            .O(N__36917),
            .I(N__36910));
    LocalMux I__7865 (
            .O(N__36914),
            .I(N__36907));
    InMux I__7864 (
            .O(N__36913),
            .I(N__36904));
    Span4Mux_h I__7863 (
            .O(N__36910),
            .I(N__36901));
    Odrv4 I__7862 (
            .O(N__36907),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__7861 (
            .O(N__36904),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__7860 (
            .O(N__36901),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__7859 (
            .O(N__36894),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__7858 (
            .O(N__36891),
            .I(N__36888));
    LocalMux I__7857 (
            .O(N__36888),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ));
    InMux I__7856 (
            .O(N__36885),
            .I(N__36881));
    InMux I__7855 (
            .O(N__36884),
            .I(N__36878));
    LocalMux I__7854 (
            .O(N__36881),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__7853 (
            .O(N__36878),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__7852 (
            .O(N__36873),
            .I(N__36870));
    LocalMux I__7851 (
            .O(N__36870),
            .I(N__36867));
    Odrv4 I__7850 (
            .O(N__36867),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ));
    InMux I__7849 (
            .O(N__36864),
            .I(N__36861));
    LocalMux I__7848 (
            .O(N__36861),
            .I(N__36857));
    InMux I__7847 (
            .O(N__36860),
            .I(N__36854));
    Odrv4 I__7846 (
            .O(N__36857),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__7845 (
            .O(N__36854),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__7844 (
            .O(N__36849),
            .I(N__36846));
    LocalMux I__7843 (
            .O(N__36846),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ));
    InMux I__7842 (
            .O(N__36843),
            .I(N__36839));
    InMux I__7841 (
            .O(N__36842),
            .I(N__36836));
    LocalMux I__7840 (
            .O(N__36839),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__7839 (
            .O(N__36836),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__7838 (
            .O(N__36831),
            .I(N__36828));
    InMux I__7837 (
            .O(N__36828),
            .I(N__36825));
    LocalMux I__7836 (
            .O(N__36825),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__7835 (
            .O(N__36822),
            .I(N__36819));
    InMux I__7834 (
            .O(N__36819),
            .I(N__36816));
    LocalMux I__7833 (
            .O(N__36816),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__7832 (
            .O(N__36813),
            .I(N__36810));
    InMux I__7831 (
            .O(N__36810),
            .I(N__36807));
    LocalMux I__7830 (
            .O(N__36807),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__7829 (
            .O(N__36804),
            .I(N__36801));
    InMux I__7828 (
            .O(N__36801),
            .I(N__36798));
    LocalMux I__7827 (
            .O(N__36798),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__7826 (
            .O(N__36795),
            .I(N__36791));
    InMux I__7825 (
            .O(N__36794),
            .I(N__36787));
    LocalMux I__7824 (
            .O(N__36791),
            .I(N__36784));
    InMux I__7823 (
            .O(N__36790),
            .I(N__36781));
    LocalMux I__7822 (
            .O(N__36787),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__7821 (
            .O(N__36784),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__7820 (
            .O(N__36781),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__7819 (
            .O(N__36774),
            .I(N__36770));
    InMux I__7818 (
            .O(N__36773),
            .I(N__36766));
    LocalMux I__7817 (
            .O(N__36770),
            .I(N__36763));
    InMux I__7816 (
            .O(N__36769),
            .I(N__36760));
    LocalMux I__7815 (
            .O(N__36766),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__7814 (
            .O(N__36763),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__7813 (
            .O(N__36760),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__7812 (
            .O(N__36753),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__7811 (
            .O(N__36750),
            .I(N__36746));
    InMux I__7810 (
            .O(N__36749),
            .I(N__36743));
    LocalMux I__7809 (
            .O(N__36746),
            .I(N__36740));
    LocalMux I__7808 (
            .O(N__36743),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__7807 (
            .O(N__36740),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__7806 (
            .O(N__36735),
            .I(N__36732));
    LocalMux I__7805 (
            .O(N__36732),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ));
    InMux I__7804 (
            .O(N__36729),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ));
    InMux I__7803 (
            .O(N__36726),
            .I(N__36722));
    InMux I__7802 (
            .O(N__36725),
            .I(N__36719));
    LocalMux I__7801 (
            .O(N__36722),
            .I(N__36716));
    LocalMux I__7800 (
            .O(N__36719),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__7799 (
            .O(N__36716),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__7798 (
            .O(N__36711),
            .I(N__36708));
    LocalMux I__7797 (
            .O(N__36708),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ));
    InMux I__7796 (
            .O(N__36705),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ));
    InMux I__7795 (
            .O(N__36702),
            .I(N__36698));
    InMux I__7794 (
            .O(N__36701),
            .I(N__36695));
    LocalMux I__7793 (
            .O(N__36698),
            .I(N__36692));
    LocalMux I__7792 (
            .O(N__36695),
            .I(N__36687));
    Span4Mux_v I__7791 (
            .O(N__36692),
            .I(N__36687));
    Odrv4 I__7790 (
            .O(N__36687),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__7789 (
            .O(N__36684),
            .I(N__36681));
    LocalMux I__7788 (
            .O(N__36681),
            .I(N__36678));
    Odrv12 I__7787 (
            .O(N__36678),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ));
    InMux I__7786 (
            .O(N__36675),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ));
    InMux I__7785 (
            .O(N__36672),
            .I(bfn_15_19_0_));
    InMux I__7784 (
            .O(N__36669),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ));
    InMux I__7783 (
            .O(N__36666),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ));
    InMux I__7782 (
            .O(N__36663),
            .I(N__36660));
    LocalMux I__7781 (
            .O(N__36660),
            .I(N__36657));
    Odrv4 I__7780 (
            .O(N__36657),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ));
    InMux I__7779 (
            .O(N__36654),
            .I(N__36651));
    LocalMux I__7778 (
            .O(N__36651),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ));
    InMux I__7777 (
            .O(N__36648),
            .I(N__36644));
    InMux I__7776 (
            .O(N__36647),
            .I(N__36641));
    LocalMux I__7775 (
            .O(N__36644),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__7774 (
            .O(N__36641),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__7773 (
            .O(N__36636),
            .I(N__36633));
    LocalMux I__7772 (
            .O(N__36633),
            .I(N__36630));
    Span4Mux_h I__7771 (
            .O(N__36630),
            .I(N__36626));
    InMux I__7770 (
            .O(N__36629),
            .I(N__36623));
    Odrv4 I__7769 (
            .O(N__36626),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__7768 (
            .O(N__36623),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__7767 (
            .O(N__36618),
            .I(N__36615));
    LocalMux I__7766 (
            .O(N__36615),
            .I(N__36612));
    Span4Mux_h I__7765 (
            .O(N__36612),
            .I(N__36609));
    Odrv4 I__7764 (
            .O(N__36609),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ));
    InMux I__7763 (
            .O(N__36606),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ));
    InMux I__7762 (
            .O(N__36603),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ));
    InMux I__7761 (
            .O(N__36600),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ));
    InMux I__7760 (
            .O(N__36597),
            .I(bfn_15_18_0_));
    InMux I__7759 (
            .O(N__36594),
            .I(N__36590));
    InMux I__7758 (
            .O(N__36593),
            .I(N__36587));
    LocalMux I__7757 (
            .O(N__36590),
            .I(N__36584));
    LocalMux I__7756 (
            .O(N__36587),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__7755 (
            .O(N__36584),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__7754 (
            .O(N__36579),
            .I(N__36576));
    LocalMux I__7753 (
            .O(N__36576),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ));
    InMux I__7752 (
            .O(N__36573),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ));
    InMux I__7751 (
            .O(N__36570),
            .I(N__36566));
    InMux I__7750 (
            .O(N__36569),
            .I(N__36563));
    LocalMux I__7749 (
            .O(N__36566),
            .I(N__36560));
    LocalMux I__7748 (
            .O(N__36563),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__7747 (
            .O(N__36560),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__7746 (
            .O(N__36555),
            .I(N__36552));
    LocalMux I__7745 (
            .O(N__36552),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ));
    InMux I__7744 (
            .O(N__36549),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ));
    InMux I__7743 (
            .O(N__36546),
            .I(N__36542));
    InMux I__7742 (
            .O(N__36545),
            .I(N__36539));
    LocalMux I__7741 (
            .O(N__36542),
            .I(N__36536));
    LocalMux I__7740 (
            .O(N__36539),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__7739 (
            .O(N__36536),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__7738 (
            .O(N__36531),
            .I(N__36528));
    LocalMux I__7737 (
            .O(N__36528),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ));
    InMux I__7736 (
            .O(N__36525),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ));
    InMux I__7735 (
            .O(N__36522),
            .I(N__36519));
    LocalMux I__7734 (
            .O(N__36519),
            .I(N__36516));
    Span4Mux_v I__7733 (
            .O(N__36516),
            .I(N__36512));
    InMux I__7732 (
            .O(N__36515),
            .I(N__36509));
    Odrv4 I__7731 (
            .O(N__36512),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__7730 (
            .O(N__36509),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__7729 (
            .O(N__36504),
            .I(N__36501));
    LocalMux I__7728 (
            .O(N__36501),
            .I(N__36498));
    Span4Mux_v I__7727 (
            .O(N__36498),
            .I(N__36495));
    Odrv4 I__7726 (
            .O(N__36495),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ));
    InMux I__7725 (
            .O(N__36492),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ));
    CascadeMux I__7724 (
            .O(N__36489),
            .I(N__36485));
    CascadeMux I__7723 (
            .O(N__36488),
            .I(N__36482));
    InMux I__7722 (
            .O(N__36485),
            .I(N__36479));
    InMux I__7721 (
            .O(N__36482),
            .I(N__36476));
    LocalMux I__7720 (
            .O(N__36479),
            .I(N__36472));
    LocalMux I__7719 (
            .O(N__36476),
            .I(N__36469));
    CascadeMux I__7718 (
            .O(N__36475),
            .I(N__36466));
    Span4Mux_h I__7717 (
            .O(N__36472),
            .I(N__36463));
    Span4Mux_h I__7716 (
            .O(N__36469),
            .I(N__36460));
    InMux I__7715 (
            .O(N__36466),
            .I(N__36457));
    Span4Mux_v I__7714 (
            .O(N__36463),
            .I(N__36454));
    Span4Mux_v I__7713 (
            .O(N__36460),
            .I(N__36451));
    LocalMux I__7712 (
            .O(N__36457),
            .I(N__36448));
    Odrv4 I__7711 (
            .O(N__36454),
            .I(measured_delay_tr_1));
    Odrv4 I__7710 (
            .O(N__36451),
            .I(measured_delay_tr_1));
    Odrv4 I__7709 (
            .O(N__36448),
            .I(measured_delay_tr_1));
    InMux I__7708 (
            .O(N__36441),
            .I(N__36435));
    InMux I__7707 (
            .O(N__36440),
            .I(N__36435));
    LocalMux I__7706 (
            .O(N__36435),
            .I(N__36427));
    InMux I__7705 (
            .O(N__36434),
            .I(N__36416));
    InMux I__7704 (
            .O(N__36433),
            .I(N__36416));
    InMux I__7703 (
            .O(N__36432),
            .I(N__36416));
    InMux I__7702 (
            .O(N__36431),
            .I(N__36416));
    InMux I__7701 (
            .O(N__36430),
            .I(N__36416));
    Span4Mux_v I__7700 (
            .O(N__36427),
            .I(N__36410));
    LocalMux I__7699 (
            .O(N__36416),
            .I(N__36410));
    InMux I__7698 (
            .O(N__36415),
            .I(N__36407));
    Odrv4 I__7697 (
            .O(N__36410),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    LocalMux I__7696 (
            .O(N__36407),
            .I(\delay_measurement_inst.un3_elapsed_time_tr_0_i ));
    CascadeMux I__7695 (
            .O(N__36402),
            .I(N__36399));
    InMux I__7694 (
            .O(N__36399),
            .I(N__36392));
    InMux I__7693 (
            .O(N__36398),
            .I(N__36392));
    CascadeMux I__7692 (
            .O(N__36397),
            .I(N__36389));
    LocalMux I__7691 (
            .O(N__36392),
            .I(N__36384));
    InMux I__7690 (
            .O(N__36389),
            .I(N__36377));
    InMux I__7689 (
            .O(N__36388),
            .I(N__36377));
    InMux I__7688 (
            .O(N__36387),
            .I(N__36377));
    Odrv12 I__7687 (
            .O(N__36384),
            .I(\delay_measurement_inst.delay_tr_reg_5_tz_1 ));
    LocalMux I__7686 (
            .O(N__36377),
            .I(\delay_measurement_inst.delay_tr_reg_5_tz_1 ));
    InMux I__7685 (
            .O(N__36372),
            .I(N__36369));
    LocalMux I__7684 (
            .O(N__36369),
            .I(N__36364));
    InMux I__7683 (
            .O(N__36368),
            .I(N__36361));
    InMux I__7682 (
            .O(N__36367),
            .I(N__36358));
    Span4Mux_v I__7681 (
            .O(N__36364),
            .I(N__36353));
    LocalMux I__7680 (
            .O(N__36361),
            .I(N__36353));
    LocalMux I__7679 (
            .O(N__36358),
            .I(N__36350));
    Span4Mux_v I__7678 (
            .O(N__36353),
            .I(N__36344));
    Span4Mux_v I__7677 (
            .O(N__36350),
            .I(N__36344));
    InMux I__7676 (
            .O(N__36349),
            .I(N__36341));
    Span4Mux_h I__7675 (
            .O(N__36344),
            .I(N__36338));
    LocalMux I__7674 (
            .O(N__36341),
            .I(measured_delay_tr_2));
    Odrv4 I__7673 (
            .O(N__36338),
            .I(measured_delay_tr_2));
    CascadeMux I__7672 (
            .O(N__36333),
            .I(N__36329));
    InMux I__7671 (
            .O(N__36332),
            .I(N__36325));
    InMux I__7670 (
            .O(N__36329),
            .I(N__36322));
    InMux I__7669 (
            .O(N__36328),
            .I(N__36319));
    LocalMux I__7668 (
            .O(N__36325),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__7667 (
            .O(N__36322),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__7666 (
            .O(N__36319),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__7665 (
            .O(N__36312),
            .I(N__36309));
    LocalMux I__7664 (
            .O(N__36309),
            .I(N__36306));
    Span4Mux_v I__7663 (
            .O(N__36306),
            .I(N__36302));
    InMux I__7662 (
            .O(N__36305),
            .I(N__36299));
    Odrv4 I__7661 (
            .O(N__36302),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__7660 (
            .O(N__36299),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__7659 (
            .O(N__36294),
            .I(N__36291));
    LocalMux I__7658 (
            .O(N__36291),
            .I(N__36288));
    Span4Mux_v I__7657 (
            .O(N__36288),
            .I(N__36285));
    Odrv4 I__7656 (
            .O(N__36285),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ));
    InMux I__7655 (
            .O(N__36282),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ));
    InMux I__7654 (
            .O(N__36279),
            .I(N__36276));
    LocalMux I__7653 (
            .O(N__36276),
            .I(N__36273));
    Span4Mux_h I__7652 (
            .O(N__36273),
            .I(N__36269));
    InMux I__7651 (
            .O(N__36272),
            .I(N__36266));
    Odrv4 I__7650 (
            .O(N__36269),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__7649 (
            .O(N__36266),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__7648 (
            .O(N__36261),
            .I(N__36258));
    InMux I__7647 (
            .O(N__36258),
            .I(N__36255));
    LocalMux I__7646 (
            .O(N__36255),
            .I(N__36252));
    Span4Mux_h I__7645 (
            .O(N__36252),
            .I(N__36249));
    Odrv4 I__7644 (
            .O(N__36249),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ));
    InMux I__7643 (
            .O(N__36246),
            .I(N__36243));
    LocalMux I__7642 (
            .O(N__36243),
            .I(N__36240));
    Span12Mux_h I__7641 (
            .O(N__36240),
            .I(N__36237));
    Odrv12 I__7640 (
            .O(N__36237),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ));
    InMux I__7639 (
            .O(N__36234),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ));
    InMux I__7638 (
            .O(N__36231),
            .I(N__36228));
    LocalMux I__7637 (
            .O(N__36228),
            .I(N__36225));
    Span4Mux_h I__7636 (
            .O(N__36225),
            .I(N__36221));
    InMux I__7635 (
            .O(N__36224),
            .I(N__36218));
    Odrv4 I__7634 (
            .O(N__36221),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__7633 (
            .O(N__36218),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__7632 (
            .O(N__36213),
            .I(N__36210));
    LocalMux I__7631 (
            .O(N__36210),
            .I(N__36207));
    Span4Mux_v I__7630 (
            .O(N__36207),
            .I(N__36204));
    Odrv4 I__7629 (
            .O(N__36204),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ));
    InMux I__7628 (
            .O(N__36201),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ));
    InMux I__7627 (
            .O(N__36198),
            .I(N__36195));
    LocalMux I__7626 (
            .O(N__36195),
            .I(N__36192));
    Span4Mux_h I__7625 (
            .O(N__36192),
            .I(N__36188));
    InMux I__7624 (
            .O(N__36191),
            .I(N__36185));
    Odrv4 I__7623 (
            .O(N__36188),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__7622 (
            .O(N__36185),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__7621 (
            .O(N__36180),
            .I(N__36177));
    LocalMux I__7620 (
            .O(N__36177),
            .I(N__36174));
    Span4Mux_h I__7619 (
            .O(N__36174),
            .I(N__36171));
    Odrv4 I__7618 (
            .O(N__36171),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ));
    InMux I__7617 (
            .O(N__36168),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ));
    InMux I__7616 (
            .O(N__36165),
            .I(N__36162));
    LocalMux I__7615 (
            .O(N__36162),
            .I(N__36159));
    Span4Mux_h I__7614 (
            .O(N__36159),
            .I(N__36156));
    Odrv4 I__7613 (
            .O(N__36156),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__7612 (
            .O(N__36153),
            .I(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0_cascade_ ));
    InMux I__7611 (
            .O(N__36150),
            .I(N__36145));
    InMux I__7610 (
            .O(N__36149),
            .I(N__36142));
    InMux I__7609 (
            .O(N__36148),
            .I(N__36139));
    LocalMux I__7608 (
            .O(N__36145),
            .I(N__36136));
    LocalMux I__7607 (
            .O(N__36142),
            .I(N__36131));
    LocalMux I__7606 (
            .O(N__36139),
            .I(N__36131));
    Span4Mux_h I__7605 (
            .O(N__36136),
            .I(N__36126));
    Span4Mux_v I__7604 (
            .O(N__36131),
            .I(N__36126));
    Span4Mux_v I__7603 (
            .O(N__36126),
            .I(N__36123));
    Span4Mux_v I__7602 (
            .O(N__36123),
            .I(N__36120));
    Odrv4 I__7601 (
            .O(N__36120),
            .I(il_max_comp1_D2));
    InMux I__7600 (
            .O(N__36117),
            .I(N__36112));
    InMux I__7599 (
            .O(N__36116),
            .I(N__36107));
    CascadeMux I__7598 (
            .O(N__36115),
            .I(N__36104));
    LocalMux I__7597 (
            .O(N__36112),
            .I(N__36101));
    InMux I__7596 (
            .O(N__36111),
            .I(N__36096));
    InMux I__7595 (
            .O(N__36110),
            .I(N__36096));
    LocalMux I__7594 (
            .O(N__36107),
            .I(N__36092));
    InMux I__7593 (
            .O(N__36104),
            .I(N__36089));
    Span4Mux_h I__7592 (
            .O(N__36101),
            .I(N__36086));
    LocalMux I__7591 (
            .O(N__36096),
            .I(N__36083));
    InMux I__7590 (
            .O(N__36095),
            .I(N__36080));
    Odrv4 I__7589 (
            .O(N__36092),
            .I(state_3));
    LocalMux I__7588 (
            .O(N__36089),
            .I(state_3));
    Odrv4 I__7587 (
            .O(N__36086),
            .I(state_3));
    Odrv4 I__7586 (
            .O(N__36083),
            .I(state_3));
    LocalMux I__7585 (
            .O(N__36080),
            .I(state_3));
    InMux I__7584 (
            .O(N__36069),
            .I(N__36066));
    LocalMux I__7583 (
            .O(N__36066),
            .I(N__36061));
    InMux I__7582 (
            .O(N__36065),
            .I(N__36058));
    InMux I__7581 (
            .O(N__36064),
            .I(N__36055));
    Odrv4 I__7580 (
            .O(N__36061),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__7579 (
            .O(N__36058),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__7578 (
            .O(N__36055),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__7577 (
            .O(N__36048),
            .I(N__36045));
    InMux I__7576 (
            .O(N__36045),
            .I(N__36041));
    CascadeMux I__7575 (
            .O(N__36044),
            .I(N__36037));
    LocalMux I__7574 (
            .O(N__36041),
            .I(N__36033));
    InMux I__7573 (
            .O(N__36040),
            .I(N__36026));
    InMux I__7572 (
            .O(N__36037),
            .I(N__36026));
    InMux I__7571 (
            .O(N__36036),
            .I(N__36026));
    Odrv12 I__7570 (
            .O(N__36033),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__7569 (
            .O(N__36026),
            .I(\phase_controller_inst1.hc_time_passed ));
    IoInMux I__7568 (
            .O(N__36021),
            .I(N__36018));
    LocalMux I__7567 (
            .O(N__36018),
            .I(N__36015));
    IoSpan4Mux I__7566 (
            .O(N__36015),
            .I(N__36012));
    Span4Mux_s2_v I__7565 (
            .O(N__36012),
            .I(N__36009));
    Sp12to4 I__7564 (
            .O(N__36009),
            .I(N__36006));
    Span12Mux_v I__7563 (
            .O(N__36006),
            .I(N__36003));
    Odrv12 I__7562 (
            .O(N__36003),
            .I(s2_phy_c));
    CascadeMux I__7561 (
            .O(N__36000),
            .I(\delay_measurement_inst.N_384_cascade_ ));
    InMux I__7560 (
            .O(N__35997),
            .I(N__35993));
    CascadeMux I__7559 (
            .O(N__35996),
            .I(N__35990));
    LocalMux I__7558 (
            .O(N__35993),
            .I(N__35986));
    InMux I__7557 (
            .O(N__35990),
            .I(N__35983));
    InMux I__7556 (
            .O(N__35989),
            .I(N__35979));
    Span4Mux_v I__7555 (
            .O(N__35986),
            .I(N__35974));
    LocalMux I__7554 (
            .O(N__35983),
            .I(N__35974));
    CascadeMux I__7553 (
            .O(N__35982),
            .I(N__35971));
    LocalMux I__7552 (
            .O(N__35979),
            .I(N__35968));
    Span4Mux_v I__7551 (
            .O(N__35974),
            .I(N__35965));
    InMux I__7550 (
            .O(N__35971),
            .I(N__35962));
    Span12Mux_v I__7549 (
            .O(N__35968),
            .I(N__35959));
    Span4Mux_v I__7548 (
            .O(N__35965),
            .I(N__35956));
    LocalMux I__7547 (
            .O(N__35962),
            .I(measured_delay_tr_4));
    Odrv12 I__7546 (
            .O(N__35959),
            .I(measured_delay_tr_4));
    Odrv4 I__7545 (
            .O(N__35956),
            .I(measured_delay_tr_4));
    InMux I__7544 (
            .O(N__35949),
            .I(N__35945));
    InMux I__7543 (
            .O(N__35948),
            .I(N__35942));
    LocalMux I__7542 (
            .O(N__35945),
            .I(N__35938));
    LocalMux I__7541 (
            .O(N__35942),
            .I(N__35935));
    InMux I__7540 (
            .O(N__35941),
            .I(N__35932));
    Span4Mux_h I__7539 (
            .O(N__35938),
            .I(N__35927));
    Span4Mux_v I__7538 (
            .O(N__35935),
            .I(N__35927));
    LocalMux I__7537 (
            .O(N__35932),
            .I(N__35923));
    Span4Mux_h I__7536 (
            .O(N__35927),
            .I(N__35920));
    InMux I__7535 (
            .O(N__35926),
            .I(N__35917));
    Span4Mux_h I__7534 (
            .O(N__35923),
            .I(N__35914));
    Odrv4 I__7533 (
            .O(N__35920),
            .I(measured_delay_tr_5));
    LocalMux I__7532 (
            .O(N__35917),
            .I(measured_delay_tr_5));
    Odrv4 I__7531 (
            .O(N__35914),
            .I(measured_delay_tr_5));
    InMux I__7530 (
            .O(N__35907),
            .I(N__35903));
    InMux I__7529 (
            .O(N__35906),
            .I(N__35900));
    LocalMux I__7528 (
            .O(N__35903),
            .I(N__35895));
    LocalMux I__7527 (
            .O(N__35900),
            .I(N__35892));
    InMux I__7526 (
            .O(N__35899),
            .I(N__35889));
    CascadeMux I__7525 (
            .O(N__35898),
            .I(N__35886));
    Span4Mux_h I__7524 (
            .O(N__35895),
            .I(N__35883));
    Span4Mux_h I__7523 (
            .O(N__35892),
            .I(N__35878));
    LocalMux I__7522 (
            .O(N__35889),
            .I(N__35878));
    InMux I__7521 (
            .O(N__35886),
            .I(N__35875));
    Span4Mux_h I__7520 (
            .O(N__35883),
            .I(N__35872));
    Span4Mux_v I__7519 (
            .O(N__35878),
            .I(N__35869));
    LocalMux I__7518 (
            .O(N__35875),
            .I(measured_delay_tr_7));
    Odrv4 I__7517 (
            .O(N__35872),
            .I(measured_delay_tr_7));
    Odrv4 I__7516 (
            .O(N__35869),
            .I(measured_delay_tr_7));
    CascadeMux I__7515 (
            .O(N__35862),
            .I(N__35859));
    InMux I__7514 (
            .O(N__35859),
            .I(N__35853));
    InMux I__7513 (
            .O(N__35858),
            .I(N__35853));
    LocalMux I__7512 (
            .O(N__35853),
            .I(N__35849));
    InMux I__7511 (
            .O(N__35852),
            .I(N__35846));
    Odrv4 I__7510 (
            .O(N__35849),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31 ));
    LocalMux I__7509 (
            .O(N__35846),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31 ));
    InMux I__7508 (
            .O(N__35841),
            .I(N__35837));
    InMux I__7507 (
            .O(N__35840),
            .I(N__35834));
    LocalMux I__7506 (
            .O(N__35837),
            .I(N__35830));
    LocalMux I__7505 (
            .O(N__35834),
            .I(N__35827));
    InMux I__7504 (
            .O(N__35833),
            .I(N__35824));
    Span4Mux_h I__7503 (
            .O(N__35830),
            .I(N__35820));
    Span4Mux_h I__7502 (
            .O(N__35827),
            .I(N__35815));
    LocalMux I__7501 (
            .O(N__35824),
            .I(N__35815));
    InMux I__7500 (
            .O(N__35823),
            .I(N__35812));
    Span4Mux_h I__7499 (
            .O(N__35820),
            .I(N__35809));
    Span4Mux_v I__7498 (
            .O(N__35815),
            .I(N__35806));
    LocalMux I__7497 (
            .O(N__35812),
            .I(measured_delay_tr_8));
    Odrv4 I__7496 (
            .O(N__35809),
            .I(measured_delay_tr_8));
    Odrv4 I__7495 (
            .O(N__35806),
            .I(measured_delay_tr_8));
    CascadeMux I__7494 (
            .O(N__35799),
            .I(N__35796));
    InMux I__7493 (
            .O(N__35796),
            .I(N__35792));
    CascadeMux I__7492 (
            .O(N__35795),
            .I(N__35789));
    LocalMux I__7491 (
            .O(N__35792),
            .I(N__35784));
    InMux I__7490 (
            .O(N__35789),
            .I(N__35781));
    InMux I__7489 (
            .O(N__35788),
            .I(N__35778));
    CascadeMux I__7488 (
            .O(N__35787),
            .I(N__35775));
    Span4Mux_h I__7487 (
            .O(N__35784),
            .I(N__35772));
    LocalMux I__7486 (
            .O(N__35781),
            .I(N__35767));
    LocalMux I__7485 (
            .O(N__35778),
            .I(N__35767));
    InMux I__7484 (
            .O(N__35775),
            .I(N__35764));
    Span4Mux_v I__7483 (
            .O(N__35772),
            .I(N__35761));
    Span4Mux_h I__7482 (
            .O(N__35767),
            .I(N__35758));
    LocalMux I__7481 (
            .O(N__35764),
            .I(measured_delay_tr_3));
    Odrv4 I__7480 (
            .O(N__35761),
            .I(measured_delay_tr_3));
    Odrv4 I__7479 (
            .O(N__35758),
            .I(measured_delay_tr_3));
    InMux I__7478 (
            .O(N__35751),
            .I(N__35748));
    LocalMux I__7477 (
            .O(N__35748),
            .I(N__35745));
    Odrv4 I__7476 (
            .O(N__35745),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ));
    InMux I__7475 (
            .O(N__35742),
            .I(N__35739));
    LocalMux I__7474 (
            .O(N__35739),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ));
    CascadeMux I__7473 (
            .O(N__35736),
            .I(\delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31_cascade_ ));
    InMux I__7472 (
            .O(N__35733),
            .I(N__35730));
    LocalMux I__7471 (
            .O(N__35730),
            .I(N__35725));
    InMux I__7470 (
            .O(N__35729),
            .I(N__35722));
    InMux I__7469 (
            .O(N__35728),
            .I(N__35719));
    Span4Mux_h I__7468 (
            .O(N__35725),
            .I(N__35716));
    LocalMux I__7467 (
            .O(N__35722),
            .I(N__35711));
    LocalMux I__7466 (
            .O(N__35719),
            .I(N__35711));
    Odrv4 I__7465 (
            .O(N__35716),
            .I(measured_delay_tr_6));
    Odrv12 I__7464 (
            .O(N__35711),
            .I(measured_delay_tr_6));
    InMux I__7463 (
            .O(N__35706),
            .I(N__35703));
    LocalMux I__7462 (
            .O(N__35703),
            .I(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0 ));
    CascadeMux I__7461 (
            .O(N__35700),
            .I(\delay_measurement_inst.N_381_cascade_ ));
    InMux I__7460 (
            .O(N__35697),
            .I(N__35694));
    LocalMux I__7459 (
            .O(N__35694),
            .I(\delay_measurement_inst.delay_tr_timer.N_376 ));
    CascadeMux I__7458 (
            .O(N__35691),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_ ));
    CascadeMux I__7457 (
            .O(N__35688),
            .I(\delay_measurement_inst.N_498_cascade_ ));
    InMux I__7456 (
            .O(N__35685),
            .I(N__35681));
    InMux I__7455 (
            .O(N__35684),
            .I(N__35678));
    LocalMux I__7454 (
            .O(N__35681),
            .I(\delay_measurement_inst.N_381 ));
    LocalMux I__7453 (
            .O(N__35678),
            .I(\delay_measurement_inst.N_381 ));
    InMux I__7452 (
            .O(N__35673),
            .I(N__35668));
    InMux I__7451 (
            .O(N__35672),
            .I(N__35663));
    InMux I__7450 (
            .O(N__35671),
            .I(N__35663));
    LocalMux I__7449 (
            .O(N__35668),
            .I(N__35660));
    LocalMux I__7448 (
            .O(N__35663),
            .I(\delay_measurement_inst.N_384 ));
    Odrv4 I__7447 (
            .O(N__35660),
            .I(\delay_measurement_inst.N_384 ));
    InMux I__7446 (
            .O(N__35655),
            .I(N__35651));
    InMux I__7445 (
            .O(N__35654),
            .I(N__35648));
    LocalMux I__7444 (
            .O(N__35651),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__7443 (
            .O(N__35648),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__7442 (
            .O(N__35643),
            .I(N__35640));
    InMux I__7441 (
            .O(N__35640),
            .I(N__35637));
    LocalMux I__7440 (
            .O(N__35637),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ));
    InMux I__7439 (
            .O(N__35634),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__7438 (
            .O(N__35631),
            .I(N__35627));
    InMux I__7437 (
            .O(N__35630),
            .I(N__35624));
    LocalMux I__7436 (
            .O(N__35627),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__7435 (
            .O(N__35624),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__7434 (
            .O(N__35619),
            .I(N__35616));
    LocalMux I__7433 (
            .O(N__35616),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ));
    InMux I__7432 (
            .O(N__35613),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__7431 (
            .O(N__35610),
            .I(N__35606));
    InMux I__7430 (
            .O(N__35609),
            .I(N__35603));
    LocalMux I__7429 (
            .O(N__35606),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__7428 (
            .O(N__35603),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__7427 (
            .O(N__35598),
            .I(N__35595));
    InMux I__7426 (
            .O(N__35595),
            .I(N__35592));
    LocalMux I__7425 (
            .O(N__35592),
            .I(N__35589));
    Odrv4 I__7424 (
            .O(N__35589),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ));
    InMux I__7423 (
            .O(N__35586),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ));
    InMux I__7422 (
            .O(N__35583),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__7421 (
            .O(N__35580),
            .I(N__35576));
    InMux I__7420 (
            .O(N__35579),
            .I(N__35573));
    LocalMux I__7419 (
            .O(N__35576),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__7418 (
            .O(N__35573),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__7417 (
            .O(N__35568),
            .I(N__35565));
    InMux I__7416 (
            .O(N__35565),
            .I(N__35562));
    LocalMux I__7415 (
            .O(N__35562),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ));
    InMux I__7414 (
            .O(N__35559),
            .I(bfn_15_10_0_));
    InMux I__7413 (
            .O(N__35556),
            .I(N__35552));
    InMux I__7412 (
            .O(N__35555),
            .I(N__35549));
    LocalMux I__7411 (
            .O(N__35552),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__7410 (
            .O(N__35549),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__7409 (
            .O(N__35544),
            .I(N__35541));
    LocalMux I__7408 (
            .O(N__35541),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ));
    InMux I__7407 (
            .O(N__35538),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__7406 (
            .O(N__35535),
            .I(N__35531));
    InMux I__7405 (
            .O(N__35534),
            .I(N__35528));
    LocalMux I__7404 (
            .O(N__35531),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__7403 (
            .O(N__35528),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__7402 (
            .O(N__35523),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ));
    CascadeMux I__7401 (
            .O(N__35520),
            .I(N__35517));
    InMux I__7400 (
            .O(N__35517),
            .I(N__35514));
    LocalMux I__7399 (
            .O(N__35514),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ));
    InMux I__7398 (
            .O(N__35511),
            .I(N__35507));
    InMux I__7397 (
            .O(N__35510),
            .I(N__35504));
    LocalMux I__7396 (
            .O(N__35507),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__7395 (
            .O(N__35504),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__7394 (
            .O(N__35499),
            .I(N__35496));
    InMux I__7393 (
            .O(N__35496),
            .I(N__35493));
    LocalMux I__7392 (
            .O(N__35493),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ));
    InMux I__7391 (
            .O(N__35490),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ));
    InMux I__7390 (
            .O(N__35487),
            .I(N__35483));
    InMux I__7389 (
            .O(N__35486),
            .I(N__35480));
    LocalMux I__7388 (
            .O(N__35483),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__7387 (
            .O(N__35480),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7386 (
            .O(N__35475),
            .I(N__35472));
    LocalMux I__7385 (
            .O(N__35472),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ));
    InMux I__7384 (
            .O(N__35469),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__7383 (
            .O(N__35466),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__7382 (
            .O(N__35463),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__7381 (
            .O(N__35460),
            .I(bfn_15_9_0_));
    InMux I__7380 (
            .O(N__35457),
            .I(N__35453));
    InMux I__7379 (
            .O(N__35456),
            .I(N__35450));
    LocalMux I__7378 (
            .O(N__35453),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__7377 (
            .O(N__35450),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__7376 (
            .O(N__35445),
            .I(N__35442));
    LocalMux I__7375 (
            .O(N__35442),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ));
    InMux I__7374 (
            .O(N__35439),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__7373 (
            .O(N__35436),
            .I(N__35432));
    InMux I__7372 (
            .O(N__35435),
            .I(N__35429));
    LocalMux I__7371 (
            .O(N__35432),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__7370 (
            .O(N__35429),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7369 (
            .O(N__35424),
            .I(N__35421));
    LocalMux I__7368 (
            .O(N__35421),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ));
    InMux I__7367 (
            .O(N__35418),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__7366 (
            .O(N__35415),
            .I(N__35411));
    InMux I__7365 (
            .O(N__35414),
            .I(N__35408));
    LocalMux I__7364 (
            .O(N__35411),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__7363 (
            .O(N__35408),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__7362 (
            .O(N__35403),
            .I(N__35400));
    LocalMux I__7361 (
            .O(N__35400),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ));
    InMux I__7360 (
            .O(N__35397),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__7359 (
            .O(N__35394),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__7358 (
            .O(N__35391),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__7357 (
            .O(N__35388),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__7356 (
            .O(N__35385),
            .I(N__35382));
    LocalMux I__7355 (
            .O(N__35382),
            .I(il_min_comp1_D1));
    CEMux I__7354 (
            .O(N__35379),
            .I(N__35375));
    CEMux I__7353 (
            .O(N__35378),
            .I(N__35371));
    LocalMux I__7352 (
            .O(N__35375),
            .I(N__35366));
    CEMux I__7351 (
            .O(N__35374),
            .I(N__35363));
    LocalMux I__7350 (
            .O(N__35371),
            .I(N__35360));
    CEMux I__7349 (
            .O(N__35370),
            .I(N__35357));
    CEMux I__7348 (
            .O(N__35369),
            .I(N__35354));
    Span4Mux_h I__7347 (
            .O(N__35366),
            .I(N__35351));
    LocalMux I__7346 (
            .O(N__35363),
            .I(N__35348));
    Span4Mux_h I__7345 (
            .O(N__35360),
            .I(N__35341));
    LocalMux I__7344 (
            .O(N__35357),
            .I(N__35341));
    LocalMux I__7343 (
            .O(N__35354),
            .I(N__35341));
    Span4Mux_h I__7342 (
            .O(N__35351),
            .I(N__35338));
    Span4Mux_h I__7341 (
            .O(N__35348),
            .I(N__35335));
    Span4Mux_v I__7340 (
            .O(N__35341),
            .I(N__35332));
    Odrv4 I__7339 (
            .O(N__35338),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__7338 (
            .O(N__35335),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__7337 (
            .O(N__35332),
            .I(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__7336 (
            .O(N__35325),
            .I(N__35322));
    LocalMux I__7335 (
            .O(N__35322),
            .I(N__35319));
    Odrv4 I__7334 (
            .O(N__35319),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ));
    CascadeMux I__7333 (
            .O(N__35316),
            .I(N__35312));
    InMux I__7332 (
            .O(N__35315),
            .I(N__35308));
    InMux I__7331 (
            .O(N__35312),
            .I(N__35305));
    InMux I__7330 (
            .O(N__35311),
            .I(N__35302));
    LocalMux I__7329 (
            .O(N__35308),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__7328 (
            .O(N__35305),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__7327 (
            .O(N__35302),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__7326 (
            .O(N__35295),
            .I(N__35291));
    InMux I__7325 (
            .O(N__35294),
            .I(N__35288));
    LocalMux I__7324 (
            .O(N__35291),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__7323 (
            .O(N__35288),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7322 (
            .O(N__35283),
            .I(N__35280));
    LocalMux I__7321 (
            .O(N__35280),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ));
    InMux I__7320 (
            .O(N__35277),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__7319 (
            .O(N__35274),
            .I(N__35271));
    LocalMux I__7318 (
            .O(N__35271),
            .I(N__35268));
    Odrv4 I__7317 (
            .O(N__35268),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ));
    CascadeMux I__7316 (
            .O(N__35265),
            .I(N__35262));
    InMux I__7315 (
            .O(N__35262),
            .I(N__35258));
    InMux I__7314 (
            .O(N__35261),
            .I(N__35255));
    LocalMux I__7313 (
            .O(N__35258),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__7312 (
            .O(N__35255),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__7311 (
            .O(N__35250),
            .I(N__35247));
    InMux I__7310 (
            .O(N__35247),
            .I(N__35244));
    LocalMux I__7309 (
            .O(N__35244),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ));
    InMux I__7308 (
            .O(N__35241),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__7307 (
            .O(N__35238),
            .I(N__35234));
    InMux I__7306 (
            .O(N__35237),
            .I(N__35231));
    LocalMux I__7305 (
            .O(N__35234),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__7304 (
            .O(N__35231),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__7303 (
            .O(N__35226),
            .I(N__35223));
    LocalMux I__7302 (
            .O(N__35223),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ));
    InMux I__7301 (
            .O(N__35220),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__7300 (
            .O(N__35217),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__7299 (
            .O(N__35214),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__7298 (
            .O(N__35211),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__7297 (
            .O(N__35208),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__7296 (
            .O(N__35205),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__7295 (
            .O(N__35202),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__7294 (
            .O(N__35199),
            .I(bfn_14_28_0_));
    InMux I__7293 (
            .O(N__35196),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__7292 (
            .O(N__35193),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__7291 (
            .O(N__35190),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__7290 (
            .O(N__35187),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__7289 (
            .O(N__35184),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__7288 (
            .O(N__35181),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__7287 (
            .O(N__35178),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__7286 (
            .O(N__35175),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__7285 (
            .O(N__35172),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__7284 (
            .O(N__35169),
            .I(bfn_14_27_0_));
    InMux I__7283 (
            .O(N__35166),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__7282 (
            .O(N__35163),
            .I(bfn_14_25_0_));
    InMux I__7281 (
            .O(N__35160),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__7280 (
            .O(N__35157),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__7279 (
            .O(N__35154),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__7278 (
            .O(N__35151),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__7277 (
            .O(N__35148),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__7276 (
            .O(N__35145),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__7275 (
            .O(N__35142),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__7274 (
            .O(N__35139),
            .I(bfn_14_26_0_));
    InMux I__7273 (
            .O(N__35136),
            .I(N__35133));
    LocalMux I__7272 (
            .O(N__35133),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ));
    InMux I__7271 (
            .O(N__35130),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__7270 (
            .O(N__35127),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ));
    CascadeMux I__7269 (
            .O(N__35124),
            .I(N__35121));
    InMux I__7268 (
            .O(N__35121),
            .I(N__35118));
    LocalMux I__7267 (
            .O(N__35118),
            .I(N__35115));
    Odrv4 I__7266 (
            .O(N__35115),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__7265 (
            .O(N__35112),
            .I(N__35109));
    LocalMux I__7264 (
            .O(N__35109),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__7263 (
            .O(N__35106),
            .I(N__35103));
    InMux I__7262 (
            .O(N__35103),
            .I(N__35100));
    LocalMux I__7261 (
            .O(N__35100),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__7260 (
            .O(N__35097),
            .I(N__35094));
    LocalMux I__7259 (
            .O(N__35094),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__7258 (
            .O(N__35091),
            .I(N__35088));
    InMux I__7257 (
            .O(N__35088),
            .I(N__35085));
    LocalMux I__7256 (
            .O(N__35085),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__7255 (
            .O(N__35082),
            .I(N__35079));
    LocalMux I__7254 (
            .O(N__35079),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__7253 (
            .O(N__35076),
            .I(N__35073));
    LocalMux I__7252 (
            .O(N__35073),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__7251 (
            .O(N__35070),
            .I(N__35067));
    LocalMux I__7250 (
            .O(N__35067),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__7249 (
            .O(N__35064),
            .I(N__35061));
    LocalMux I__7248 (
            .O(N__35061),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ));
    InMux I__7247 (
            .O(N__35058),
            .I(N__35055));
    LocalMux I__7246 (
            .O(N__35055),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ));
    InMux I__7245 (
            .O(N__35052),
            .I(N__35049));
    LocalMux I__7244 (
            .O(N__35049),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ));
    InMux I__7243 (
            .O(N__35046),
            .I(N__35043));
    LocalMux I__7242 (
            .O(N__35043),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    CascadeMux I__7241 (
            .O(N__35040),
            .I(N__35037));
    InMux I__7240 (
            .O(N__35037),
            .I(N__35034));
    LocalMux I__7239 (
            .O(N__35034),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__7238 (
            .O(N__35031),
            .I(N__35028));
    LocalMux I__7237 (
            .O(N__35028),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__7236 (
            .O(N__35025),
            .I(N__35022));
    LocalMux I__7235 (
            .O(N__35022),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__7234 (
            .O(N__35019),
            .I(N__35016));
    LocalMux I__7233 (
            .O(N__35016),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__7232 (
            .O(N__35013),
            .I(N__35010));
    LocalMux I__7231 (
            .O(N__35010),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__7230 (
            .O(N__35007),
            .I(N__35004));
    LocalMux I__7229 (
            .O(N__35004),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__7228 (
            .O(N__35001),
            .I(N__34998));
    InMux I__7227 (
            .O(N__34998),
            .I(N__34995));
    LocalMux I__7226 (
            .O(N__34995),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__7225 (
            .O(N__34992),
            .I(N__34989));
    InMux I__7224 (
            .O(N__34989),
            .I(N__34986));
    LocalMux I__7223 (
            .O(N__34986),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__7222 (
            .O(N__34983),
            .I(N__34980));
    LocalMux I__7221 (
            .O(N__34980),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__7220 (
            .O(N__34977),
            .I(N__34974));
    InMux I__7219 (
            .O(N__34974),
            .I(N__34971));
    LocalMux I__7218 (
            .O(N__34971),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__7217 (
            .O(N__34968),
            .I(N__34965));
    LocalMux I__7216 (
            .O(N__34965),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__7215 (
            .O(N__34962),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__7214 (
            .O(N__34959),
            .I(N__34956));
    LocalMux I__7213 (
            .O(N__34956),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ));
    CascadeMux I__7212 (
            .O(N__34953),
            .I(N__34950));
    InMux I__7211 (
            .O(N__34950),
            .I(N__34947));
    LocalMux I__7210 (
            .O(N__34947),
            .I(N__34944));
    Odrv4 I__7209 (
            .O(N__34944),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__7208 (
            .O(N__34941),
            .I(N__34938));
    LocalMux I__7207 (
            .O(N__34938),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__7206 (
            .O(N__34935),
            .I(N__34932));
    LocalMux I__7205 (
            .O(N__34932),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__7204 (
            .O(N__34929),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__7203 (
            .O(N__34926),
            .I(N__34923));
    InMux I__7202 (
            .O(N__34923),
            .I(N__34919));
    InMux I__7201 (
            .O(N__34922),
            .I(N__34916));
    LocalMux I__7200 (
            .O(N__34919),
            .I(N__34910));
    LocalMux I__7199 (
            .O(N__34916),
            .I(N__34910));
    InMux I__7198 (
            .O(N__34915),
            .I(N__34907));
    Span4Mux_v I__7197 (
            .O(N__34910),
            .I(N__34904));
    LocalMux I__7196 (
            .O(N__34907),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__7195 (
            .O(N__34904),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__7194 (
            .O(N__34899),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__7193 (
            .O(N__34896),
            .I(N__34889));
    InMux I__7192 (
            .O(N__34895),
            .I(N__34889));
    InMux I__7191 (
            .O(N__34894),
            .I(N__34886));
    LocalMux I__7190 (
            .O(N__34889),
            .I(N__34883));
    LocalMux I__7189 (
            .O(N__34886),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__7188 (
            .O(N__34883),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__7187 (
            .O(N__34878),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__7186 (
            .O(N__34875),
            .I(N__34871));
    InMux I__7185 (
            .O(N__34874),
            .I(N__34868));
    LocalMux I__7184 (
            .O(N__34871),
            .I(N__34865));
    LocalMux I__7183 (
            .O(N__34868),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__7182 (
            .O(N__34865),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__7181 (
            .O(N__34860),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__7180 (
            .O(N__34857),
            .I(N__34821));
    InMux I__7179 (
            .O(N__34856),
            .I(N__34821));
    InMux I__7178 (
            .O(N__34855),
            .I(N__34821));
    InMux I__7177 (
            .O(N__34854),
            .I(N__34821));
    InMux I__7176 (
            .O(N__34853),
            .I(N__34812));
    InMux I__7175 (
            .O(N__34852),
            .I(N__34812));
    InMux I__7174 (
            .O(N__34851),
            .I(N__34812));
    InMux I__7173 (
            .O(N__34850),
            .I(N__34812));
    InMux I__7172 (
            .O(N__34849),
            .I(N__34803));
    InMux I__7171 (
            .O(N__34848),
            .I(N__34803));
    InMux I__7170 (
            .O(N__34847),
            .I(N__34803));
    InMux I__7169 (
            .O(N__34846),
            .I(N__34803));
    InMux I__7168 (
            .O(N__34845),
            .I(N__34794));
    InMux I__7167 (
            .O(N__34844),
            .I(N__34794));
    InMux I__7166 (
            .O(N__34843),
            .I(N__34794));
    InMux I__7165 (
            .O(N__34842),
            .I(N__34794));
    InMux I__7164 (
            .O(N__34841),
            .I(N__34785));
    InMux I__7163 (
            .O(N__34840),
            .I(N__34785));
    InMux I__7162 (
            .O(N__34839),
            .I(N__34785));
    InMux I__7161 (
            .O(N__34838),
            .I(N__34785));
    InMux I__7160 (
            .O(N__34837),
            .I(N__34776));
    InMux I__7159 (
            .O(N__34836),
            .I(N__34776));
    InMux I__7158 (
            .O(N__34835),
            .I(N__34776));
    InMux I__7157 (
            .O(N__34834),
            .I(N__34776));
    InMux I__7156 (
            .O(N__34833),
            .I(N__34765));
    InMux I__7155 (
            .O(N__34832),
            .I(N__34765));
    InMux I__7154 (
            .O(N__34831),
            .I(N__34765));
    InMux I__7153 (
            .O(N__34830),
            .I(N__34765));
    LocalMux I__7152 (
            .O(N__34821),
            .I(N__34760));
    LocalMux I__7151 (
            .O(N__34812),
            .I(N__34760));
    LocalMux I__7150 (
            .O(N__34803),
            .I(N__34751));
    LocalMux I__7149 (
            .O(N__34794),
            .I(N__34751));
    LocalMux I__7148 (
            .O(N__34785),
            .I(N__34751));
    LocalMux I__7147 (
            .O(N__34776),
            .I(N__34751));
    InMux I__7146 (
            .O(N__34775),
            .I(N__34746));
    InMux I__7145 (
            .O(N__34774),
            .I(N__34746));
    LocalMux I__7144 (
            .O(N__34765),
            .I(N__34739));
    Span4Mux_v I__7143 (
            .O(N__34760),
            .I(N__34739));
    Span4Mux_v I__7142 (
            .O(N__34751),
            .I(N__34739));
    LocalMux I__7141 (
            .O(N__34746),
            .I(N__34736));
    Span4Mux_v I__7140 (
            .O(N__34739),
            .I(N__34733));
    Span4Mux_h I__7139 (
            .O(N__34736),
            .I(N__34730));
    Span4Mux_h I__7138 (
            .O(N__34733),
            .I(N__34727));
    Odrv4 I__7137 (
            .O(N__34730),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__7136 (
            .O(N__34727),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__7135 (
            .O(N__34722),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__7134 (
            .O(N__34719),
            .I(N__34716));
    InMux I__7133 (
            .O(N__34716),
            .I(N__34712));
    InMux I__7132 (
            .O(N__34715),
            .I(N__34709));
    LocalMux I__7131 (
            .O(N__34712),
            .I(N__34706));
    LocalMux I__7130 (
            .O(N__34709),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__7129 (
            .O(N__34706),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__7128 (
            .O(N__34701),
            .I(N__34697));
    CEMux I__7127 (
            .O(N__34700),
            .I(N__34692));
    LocalMux I__7126 (
            .O(N__34697),
            .I(N__34689));
    CEMux I__7125 (
            .O(N__34696),
            .I(N__34686));
    CEMux I__7124 (
            .O(N__34695),
            .I(N__34683));
    LocalMux I__7123 (
            .O(N__34692),
            .I(N__34680));
    Span4Mux_v I__7122 (
            .O(N__34689),
            .I(N__34675));
    LocalMux I__7121 (
            .O(N__34686),
            .I(N__34675));
    LocalMux I__7120 (
            .O(N__34683),
            .I(N__34672));
    Span4Mux_v I__7119 (
            .O(N__34680),
            .I(N__34667));
    Span4Mux_h I__7118 (
            .O(N__34675),
            .I(N__34667));
    Span4Mux_h I__7117 (
            .O(N__34672),
            .I(N__34664));
    Span4Mux_v I__7116 (
            .O(N__34667),
            .I(N__34661));
    Span4Mux_h I__7115 (
            .O(N__34664),
            .I(N__34658));
    Odrv4 I__7114 (
            .O(N__34661),
            .I(\current_shift_inst.timer_s1.N_186_i ));
    Odrv4 I__7113 (
            .O(N__34658),
            .I(\current_shift_inst.timer_s1.N_186_i ));
    InMux I__7112 (
            .O(N__34653),
            .I(N__34649));
    InMux I__7111 (
            .O(N__34652),
            .I(N__34646));
    LocalMux I__7110 (
            .O(N__34649),
            .I(N__34643));
    LocalMux I__7109 (
            .O(N__34646),
            .I(N__34640));
    Span4Mux_v I__7108 (
            .O(N__34643),
            .I(N__34637));
    Span4Mux_h I__7107 (
            .O(N__34640),
            .I(N__34634));
    Odrv4 I__7106 (
            .O(N__34637),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__7105 (
            .O(N__34634),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__7104 (
            .O(N__34629),
            .I(N__34626));
    LocalMux I__7103 (
            .O(N__34626),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__7102 (
            .O(N__34623),
            .I(N__34620));
    InMux I__7101 (
            .O(N__34620),
            .I(N__34615));
    InMux I__7100 (
            .O(N__34619),
            .I(N__34610));
    InMux I__7099 (
            .O(N__34618),
            .I(N__34610));
    LocalMux I__7098 (
            .O(N__34615),
            .I(N__34607));
    LocalMux I__7097 (
            .O(N__34610),
            .I(N__34604));
    Span4Mux_h I__7096 (
            .O(N__34607),
            .I(N__34601));
    Span4Mux_h I__7095 (
            .O(N__34604),
            .I(N__34598));
    Span4Mux_h I__7094 (
            .O(N__34601),
            .I(N__34593));
    Span4Mux_h I__7093 (
            .O(N__34598),
            .I(N__34593));
    Odrv4 I__7092 (
            .O(N__34593),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__7091 (
            .O(N__34590),
            .I(N__34553));
    CascadeMux I__7090 (
            .O(N__34589),
            .I(N__34550));
    CascadeMux I__7089 (
            .O(N__34588),
            .I(N__34547));
    CascadeMux I__7088 (
            .O(N__34587),
            .I(N__34544));
    CascadeMux I__7087 (
            .O(N__34586),
            .I(N__34541));
    CascadeMux I__7086 (
            .O(N__34585),
            .I(N__34538));
    CascadeMux I__7085 (
            .O(N__34584),
            .I(N__34535));
    CascadeMux I__7084 (
            .O(N__34583),
            .I(N__34532));
    CascadeMux I__7083 (
            .O(N__34582),
            .I(N__34529));
    CascadeMux I__7082 (
            .O(N__34581),
            .I(N__34526));
    CascadeMux I__7081 (
            .O(N__34580),
            .I(N__34523));
    CascadeMux I__7080 (
            .O(N__34579),
            .I(N__34520));
    CascadeMux I__7079 (
            .O(N__34578),
            .I(N__34517));
    CascadeMux I__7078 (
            .O(N__34577),
            .I(N__34514));
    CascadeMux I__7077 (
            .O(N__34576),
            .I(N__34511));
    InMux I__7076 (
            .O(N__34575),
            .I(N__34506));
    InMux I__7075 (
            .O(N__34574),
            .I(N__34506));
    CascadeMux I__7074 (
            .O(N__34573),
            .I(N__34503));
    CascadeMux I__7073 (
            .O(N__34572),
            .I(N__34500));
    CascadeMux I__7072 (
            .O(N__34571),
            .I(N__34497));
    CascadeMux I__7071 (
            .O(N__34570),
            .I(N__34494));
    CascadeMux I__7070 (
            .O(N__34569),
            .I(N__34491));
    CascadeMux I__7069 (
            .O(N__34568),
            .I(N__34487));
    CascadeMux I__7068 (
            .O(N__34567),
            .I(N__34484));
    InMux I__7067 (
            .O(N__34566),
            .I(N__34475));
    InMux I__7066 (
            .O(N__34565),
            .I(N__34472));
    InMux I__7065 (
            .O(N__34564),
            .I(N__34465));
    InMux I__7064 (
            .O(N__34563),
            .I(N__34465));
    InMux I__7063 (
            .O(N__34562),
            .I(N__34465));
    InMux I__7062 (
            .O(N__34561),
            .I(N__34456));
    InMux I__7061 (
            .O(N__34560),
            .I(N__34456));
    InMux I__7060 (
            .O(N__34559),
            .I(N__34456));
    InMux I__7059 (
            .O(N__34558),
            .I(N__34456));
    CascadeMux I__7058 (
            .O(N__34557),
            .I(N__34453));
    CascadeMux I__7057 (
            .O(N__34556),
            .I(N__34450));
    InMux I__7056 (
            .O(N__34553),
            .I(N__34442));
    InMux I__7055 (
            .O(N__34550),
            .I(N__34442));
    InMux I__7054 (
            .O(N__34547),
            .I(N__34442));
    InMux I__7053 (
            .O(N__34544),
            .I(N__34433));
    InMux I__7052 (
            .O(N__34541),
            .I(N__34433));
    InMux I__7051 (
            .O(N__34538),
            .I(N__34433));
    InMux I__7050 (
            .O(N__34535),
            .I(N__34433));
    InMux I__7049 (
            .O(N__34532),
            .I(N__34424));
    InMux I__7048 (
            .O(N__34529),
            .I(N__34424));
    InMux I__7047 (
            .O(N__34526),
            .I(N__34424));
    InMux I__7046 (
            .O(N__34523),
            .I(N__34424));
    InMux I__7045 (
            .O(N__34520),
            .I(N__34415));
    InMux I__7044 (
            .O(N__34517),
            .I(N__34415));
    InMux I__7043 (
            .O(N__34514),
            .I(N__34415));
    InMux I__7042 (
            .O(N__34511),
            .I(N__34415));
    LocalMux I__7041 (
            .O(N__34506),
            .I(N__34412));
    InMux I__7040 (
            .O(N__34503),
            .I(N__34405));
    InMux I__7039 (
            .O(N__34500),
            .I(N__34405));
    InMux I__7038 (
            .O(N__34497),
            .I(N__34405));
    InMux I__7037 (
            .O(N__34494),
            .I(N__34394));
    InMux I__7036 (
            .O(N__34491),
            .I(N__34394));
    InMux I__7035 (
            .O(N__34490),
            .I(N__34394));
    InMux I__7034 (
            .O(N__34487),
            .I(N__34394));
    InMux I__7033 (
            .O(N__34484),
            .I(N__34394));
    CascadeMux I__7032 (
            .O(N__34483),
            .I(N__34391));
    CascadeMux I__7031 (
            .O(N__34482),
            .I(N__34388));
    CascadeMux I__7030 (
            .O(N__34481),
            .I(N__34385));
    CascadeMux I__7029 (
            .O(N__34480),
            .I(N__34382));
    CascadeMux I__7028 (
            .O(N__34479),
            .I(N__34379));
    CascadeMux I__7027 (
            .O(N__34478),
            .I(N__34376));
    LocalMux I__7026 (
            .O(N__34475),
            .I(N__34364));
    LocalMux I__7025 (
            .O(N__34472),
            .I(N__34361));
    LocalMux I__7024 (
            .O(N__34465),
            .I(N__34356));
    LocalMux I__7023 (
            .O(N__34456),
            .I(N__34356));
    InMux I__7022 (
            .O(N__34453),
            .I(N__34353));
    InMux I__7021 (
            .O(N__34450),
            .I(N__34348));
    InMux I__7020 (
            .O(N__34449),
            .I(N__34348));
    LocalMux I__7019 (
            .O(N__34442),
            .I(N__34343));
    LocalMux I__7018 (
            .O(N__34433),
            .I(N__34343));
    LocalMux I__7017 (
            .O(N__34424),
            .I(N__34338));
    LocalMux I__7016 (
            .O(N__34415),
            .I(N__34338));
    Span4Mux_h I__7015 (
            .O(N__34412),
            .I(N__34331));
    LocalMux I__7014 (
            .O(N__34405),
            .I(N__34331));
    LocalMux I__7013 (
            .O(N__34394),
            .I(N__34331));
    InMux I__7012 (
            .O(N__34391),
            .I(N__34324));
    InMux I__7011 (
            .O(N__34388),
            .I(N__34324));
    InMux I__7010 (
            .O(N__34385),
            .I(N__34324));
    InMux I__7009 (
            .O(N__34382),
            .I(N__34315));
    InMux I__7008 (
            .O(N__34379),
            .I(N__34315));
    InMux I__7007 (
            .O(N__34376),
            .I(N__34315));
    InMux I__7006 (
            .O(N__34375),
            .I(N__34315));
    InMux I__7005 (
            .O(N__34374),
            .I(N__34312));
    InMux I__7004 (
            .O(N__34373),
            .I(N__34305));
    InMux I__7003 (
            .O(N__34372),
            .I(N__34305));
    InMux I__7002 (
            .O(N__34371),
            .I(N__34305));
    InMux I__7001 (
            .O(N__34370),
            .I(N__34296));
    InMux I__7000 (
            .O(N__34369),
            .I(N__34296));
    InMux I__6999 (
            .O(N__34368),
            .I(N__34296));
    InMux I__6998 (
            .O(N__34367),
            .I(N__34296));
    Span4Mux_s2_v I__6997 (
            .O(N__34364),
            .I(N__34293));
    Span4Mux_v I__6996 (
            .O(N__34361),
            .I(N__34287));
    Span4Mux_v I__6995 (
            .O(N__34356),
            .I(N__34280));
    LocalMux I__6994 (
            .O(N__34353),
            .I(N__34280));
    LocalMux I__6993 (
            .O(N__34348),
            .I(N__34280));
    Span4Mux_v I__6992 (
            .O(N__34343),
            .I(N__34269));
    Span4Mux_v I__6991 (
            .O(N__34338),
            .I(N__34269));
    Span4Mux_h I__6990 (
            .O(N__34331),
            .I(N__34269));
    LocalMux I__6989 (
            .O(N__34324),
            .I(N__34269));
    LocalMux I__6988 (
            .O(N__34315),
            .I(N__34269));
    LocalMux I__6987 (
            .O(N__34312),
            .I(N__34262));
    LocalMux I__6986 (
            .O(N__34305),
            .I(N__34262));
    LocalMux I__6985 (
            .O(N__34296),
            .I(N__34262));
    Span4Mux_v I__6984 (
            .O(N__34293),
            .I(N__34259));
    InMux I__6983 (
            .O(N__34292),
            .I(N__34256));
    InMux I__6982 (
            .O(N__34291),
            .I(N__34253));
    InMux I__6981 (
            .O(N__34290),
            .I(N__34250));
    Span4Mux_h I__6980 (
            .O(N__34287),
            .I(N__34245));
    Span4Mux_h I__6979 (
            .O(N__34280),
            .I(N__34245));
    Span4Mux_v I__6978 (
            .O(N__34269),
            .I(N__34242));
    Span12Mux_s11_v I__6977 (
            .O(N__34262),
            .I(N__34239));
    Sp12to4 I__6976 (
            .O(N__34259),
            .I(N__34236));
    LocalMux I__6975 (
            .O(N__34256),
            .I(N__34229));
    LocalMux I__6974 (
            .O(N__34253),
            .I(N__34229));
    LocalMux I__6973 (
            .O(N__34250),
            .I(N__34229));
    Sp12to4 I__6972 (
            .O(N__34245),
            .I(N__34226));
    Span4Mux_h I__6971 (
            .O(N__34242),
            .I(N__34223));
    Span12Mux_v I__6970 (
            .O(N__34239),
            .I(N__34216));
    Span12Mux_h I__6969 (
            .O(N__34236),
            .I(N__34216));
    Span12Mux_s6_v I__6968 (
            .O(N__34229),
            .I(N__34216));
    Odrv12 I__6967 (
            .O(N__34226),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6966 (
            .O(N__34223),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6965 (
            .O(N__34216),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__6964 (
            .O(N__34209),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    InMux I__6963 (
            .O(N__34206),
            .I(N__34202));
    InMux I__6962 (
            .O(N__34205),
            .I(N__34199));
    LocalMux I__6961 (
            .O(N__34202),
            .I(N__34196));
    LocalMux I__6960 (
            .O(N__34199),
            .I(N__34193));
    Span4Mux_h I__6959 (
            .O(N__34196),
            .I(N__34190));
    Span4Mux_v I__6958 (
            .O(N__34193),
            .I(N__34187));
    Span4Mux_v I__6957 (
            .O(N__34190),
            .I(N__34184));
    Odrv4 I__6956 (
            .O(N__34187),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__6955 (
            .O(N__34184),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__6954 (
            .O(N__34179),
            .I(N__34175));
    CascadeMux I__6953 (
            .O(N__34178),
            .I(N__34172));
    InMux I__6952 (
            .O(N__34175),
            .I(N__34169));
    InMux I__6951 (
            .O(N__34172),
            .I(N__34166));
    LocalMux I__6950 (
            .O(N__34169),
            .I(N__34161));
    LocalMux I__6949 (
            .O(N__34166),
            .I(N__34161));
    Span4Mux_h I__6948 (
            .O(N__34161),
            .I(N__34158));
    Span4Mux_h I__6947 (
            .O(N__34158),
            .I(N__34155));
    Odrv4 I__6946 (
            .O(N__34155),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__6945 (
            .O(N__34152),
            .I(N__34149));
    InMux I__6944 (
            .O(N__34149),
            .I(N__34146));
    LocalMux I__6943 (
            .O(N__34146),
            .I(N__34141));
    CascadeMux I__6942 (
            .O(N__34145),
            .I(N__34138));
    InMux I__6941 (
            .O(N__34144),
            .I(N__34135));
    Span4Mux_h I__6940 (
            .O(N__34141),
            .I(N__34132));
    InMux I__6939 (
            .O(N__34138),
            .I(N__34129));
    LocalMux I__6938 (
            .O(N__34135),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__6937 (
            .O(N__34132),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    LocalMux I__6936 (
            .O(N__34129),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__6935 (
            .O(N__34122),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__6934 (
            .O(N__34119),
            .I(N__34113));
    InMux I__6933 (
            .O(N__34118),
            .I(N__34113));
    LocalMux I__6932 (
            .O(N__34113),
            .I(N__34109));
    InMux I__6931 (
            .O(N__34112),
            .I(N__34106));
    Span4Mux_v I__6930 (
            .O(N__34109),
            .I(N__34103));
    LocalMux I__6929 (
            .O(N__34106),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__6928 (
            .O(N__34103),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__6927 (
            .O(N__34098),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__6926 (
            .O(N__34095),
            .I(N__34088));
    InMux I__6925 (
            .O(N__34094),
            .I(N__34088));
    InMux I__6924 (
            .O(N__34093),
            .I(N__34085));
    LocalMux I__6923 (
            .O(N__34088),
            .I(N__34082));
    LocalMux I__6922 (
            .O(N__34085),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__6921 (
            .O(N__34082),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__6920 (
            .O(N__34077),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__6919 (
            .O(N__34074),
            .I(N__34070));
    CascadeMux I__6918 (
            .O(N__34073),
            .I(N__34067));
    InMux I__6917 (
            .O(N__34070),
            .I(N__34062));
    InMux I__6916 (
            .O(N__34067),
            .I(N__34062));
    LocalMux I__6915 (
            .O(N__34062),
            .I(N__34058));
    InMux I__6914 (
            .O(N__34061),
            .I(N__34055));
    Span4Mux_h I__6913 (
            .O(N__34058),
            .I(N__34052));
    LocalMux I__6912 (
            .O(N__34055),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__6911 (
            .O(N__34052),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__6910 (
            .O(N__34047),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__6909 (
            .O(N__34044),
            .I(N__34040));
    CascadeMux I__6908 (
            .O(N__34043),
            .I(N__34037));
    InMux I__6907 (
            .O(N__34040),
            .I(N__34031));
    InMux I__6906 (
            .O(N__34037),
            .I(N__34031));
    InMux I__6905 (
            .O(N__34036),
            .I(N__34028));
    LocalMux I__6904 (
            .O(N__34031),
            .I(N__34025));
    LocalMux I__6903 (
            .O(N__34028),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__6902 (
            .O(N__34025),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__6901 (
            .O(N__34020),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__6900 (
            .O(N__34017),
            .I(N__34010));
    InMux I__6899 (
            .O(N__34016),
            .I(N__34010));
    InMux I__6898 (
            .O(N__34015),
            .I(N__34007));
    LocalMux I__6897 (
            .O(N__34010),
            .I(N__34004));
    LocalMux I__6896 (
            .O(N__34007),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__6895 (
            .O(N__34004),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__6894 (
            .O(N__33999),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__6893 (
            .O(N__33996),
            .I(N__33992));
    InMux I__6892 (
            .O(N__33995),
            .I(N__33989));
    InMux I__6891 (
            .O(N__33992),
            .I(N__33985));
    LocalMux I__6890 (
            .O(N__33989),
            .I(N__33982));
    InMux I__6889 (
            .O(N__33988),
            .I(N__33979));
    LocalMux I__6888 (
            .O(N__33985),
            .I(N__33974));
    Span4Mux_h I__6887 (
            .O(N__33982),
            .I(N__33974));
    LocalMux I__6886 (
            .O(N__33979),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__6885 (
            .O(N__33974),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__6884 (
            .O(N__33969),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__6883 (
            .O(N__33966),
            .I(N__33963));
    InMux I__6882 (
            .O(N__33963),
            .I(N__33958));
    CascadeMux I__6881 (
            .O(N__33962),
            .I(N__33955));
    InMux I__6880 (
            .O(N__33961),
            .I(N__33952));
    LocalMux I__6879 (
            .O(N__33958),
            .I(N__33949));
    InMux I__6878 (
            .O(N__33955),
            .I(N__33946));
    LocalMux I__6877 (
            .O(N__33952),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__6876 (
            .O(N__33949),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__6875 (
            .O(N__33946),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__6874 (
            .O(N__33939),
            .I(bfn_14_16_0_));
    CascadeMux I__6873 (
            .O(N__33936),
            .I(N__33933));
    InMux I__6872 (
            .O(N__33933),
            .I(N__33930));
    LocalMux I__6871 (
            .O(N__33930),
            .I(N__33926));
    InMux I__6870 (
            .O(N__33929),
            .I(N__33922));
    Span4Mux_v I__6869 (
            .O(N__33926),
            .I(N__33919));
    InMux I__6868 (
            .O(N__33925),
            .I(N__33916));
    LocalMux I__6867 (
            .O(N__33922),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__6866 (
            .O(N__33919),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__6865 (
            .O(N__33916),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    CascadeMux I__6864 (
            .O(N__33909),
            .I(N__33906));
    InMux I__6863 (
            .O(N__33906),
            .I(N__33903));
    LocalMux I__6862 (
            .O(N__33903),
            .I(N__33898));
    CascadeMux I__6861 (
            .O(N__33902),
            .I(N__33895));
    InMux I__6860 (
            .O(N__33901),
            .I(N__33892));
    Span4Mux_h I__6859 (
            .O(N__33898),
            .I(N__33889));
    InMux I__6858 (
            .O(N__33895),
            .I(N__33886));
    LocalMux I__6857 (
            .O(N__33892),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__6856 (
            .O(N__33889),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__6855 (
            .O(N__33886),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__6854 (
            .O(N__33879),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__6853 (
            .O(N__33876),
            .I(N__33873));
    InMux I__6852 (
            .O(N__33873),
            .I(N__33869));
    InMux I__6851 (
            .O(N__33872),
            .I(N__33866));
    LocalMux I__6850 (
            .O(N__33869),
            .I(N__33860));
    LocalMux I__6849 (
            .O(N__33866),
            .I(N__33860));
    InMux I__6848 (
            .O(N__33865),
            .I(N__33857));
    Span4Mux_v I__6847 (
            .O(N__33860),
            .I(N__33854));
    LocalMux I__6846 (
            .O(N__33857),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__6845 (
            .O(N__33854),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__6844 (
            .O(N__33849),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__6843 (
            .O(N__33846),
            .I(N__33839));
    InMux I__6842 (
            .O(N__33845),
            .I(N__33839));
    InMux I__6841 (
            .O(N__33844),
            .I(N__33836));
    LocalMux I__6840 (
            .O(N__33839),
            .I(N__33833));
    LocalMux I__6839 (
            .O(N__33836),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__6838 (
            .O(N__33833),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__6837 (
            .O(N__33828),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__6836 (
            .O(N__33825),
            .I(N__33818));
    InMux I__6835 (
            .O(N__33824),
            .I(N__33818));
    InMux I__6834 (
            .O(N__33823),
            .I(N__33815));
    LocalMux I__6833 (
            .O(N__33818),
            .I(N__33812));
    LocalMux I__6832 (
            .O(N__33815),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__6831 (
            .O(N__33812),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__6830 (
            .O(N__33807),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__6829 (
            .O(N__33804),
            .I(N__33800));
    CascadeMux I__6828 (
            .O(N__33803),
            .I(N__33797));
    InMux I__6827 (
            .O(N__33800),
            .I(N__33791));
    InMux I__6826 (
            .O(N__33797),
            .I(N__33791));
    InMux I__6825 (
            .O(N__33796),
            .I(N__33788));
    LocalMux I__6824 (
            .O(N__33791),
            .I(N__33785));
    LocalMux I__6823 (
            .O(N__33788),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__6822 (
            .O(N__33785),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__6821 (
            .O(N__33780),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__6820 (
            .O(N__33777),
            .I(N__33773));
    CascadeMux I__6819 (
            .O(N__33776),
            .I(N__33770));
    InMux I__6818 (
            .O(N__33773),
            .I(N__33765));
    InMux I__6817 (
            .O(N__33770),
            .I(N__33765));
    LocalMux I__6816 (
            .O(N__33765),
            .I(N__33761));
    InMux I__6815 (
            .O(N__33764),
            .I(N__33758));
    Span4Mux_h I__6814 (
            .O(N__33761),
            .I(N__33755));
    LocalMux I__6813 (
            .O(N__33758),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__6812 (
            .O(N__33755),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__6811 (
            .O(N__33750),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__6810 (
            .O(N__33747),
            .I(N__33741));
    InMux I__6809 (
            .O(N__33746),
            .I(N__33741));
    LocalMux I__6808 (
            .O(N__33741),
            .I(N__33737));
    InMux I__6807 (
            .O(N__33740),
            .I(N__33734));
    Span4Mux_h I__6806 (
            .O(N__33737),
            .I(N__33731));
    LocalMux I__6805 (
            .O(N__33734),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__6804 (
            .O(N__33731),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__6803 (
            .O(N__33726),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__6802 (
            .O(N__33723),
            .I(N__33720));
    InMux I__6801 (
            .O(N__33720),
            .I(N__33716));
    InMux I__6800 (
            .O(N__33719),
            .I(N__33712));
    LocalMux I__6799 (
            .O(N__33716),
            .I(N__33709));
    InMux I__6798 (
            .O(N__33715),
            .I(N__33706));
    LocalMux I__6797 (
            .O(N__33712),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__6796 (
            .O(N__33709),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__6795 (
            .O(N__33706),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__6794 (
            .O(N__33699),
            .I(bfn_14_15_0_));
    InMux I__6793 (
            .O(N__33696),
            .I(N__33692));
    InMux I__6792 (
            .O(N__33695),
            .I(N__33689));
    LocalMux I__6791 (
            .O(N__33692),
            .I(N__33685));
    LocalMux I__6790 (
            .O(N__33689),
            .I(N__33682));
    InMux I__6789 (
            .O(N__33688),
            .I(N__33679));
    Span4Mux_h I__6788 (
            .O(N__33685),
            .I(N__33676));
    Odrv12 I__6787 (
            .O(N__33682),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__6786 (
            .O(N__33679),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__6785 (
            .O(N__33676),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__6784 (
            .O(N__33669),
            .I(bfn_14_13_0_));
    InMux I__6783 (
            .O(N__33666),
            .I(N__33662));
    CascadeMux I__6782 (
            .O(N__33665),
            .I(N__33659));
    LocalMux I__6781 (
            .O(N__33662),
            .I(N__33656));
    InMux I__6780 (
            .O(N__33659),
            .I(N__33653));
    Span4Mux_v I__6779 (
            .O(N__33656),
            .I(N__33647));
    LocalMux I__6778 (
            .O(N__33653),
            .I(N__33647));
    InMux I__6777 (
            .O(N__33652),
            .I(N__33644));
    Span4Mux_h I__6776 (
            .O(N__33647),
            .I(N__33641));
    LocalMux I__6775 (
            .O(N__33644),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__6774 (
            .O(N__33641),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__6773 (
            .O(N__33636),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__6772 (
            .O(N__33633),
            .I(N__33629));
    CascadeMux I__6771 (
            .O(N__33632),
            .I(N__33626));
    InMux I__6770 (
            .O(N__33629),
            .I(N__33620));
    InMux I__6769 (
            .O(N__33626),
            .I(N__33620));
    InMux I__6768 (
            .O(N__33625),
            .I(N__33617));
    LocalMux I__6767 (
            .O(N__33620),
            .I(N__33614));
    LocalMux I__6766 (
            .O(N__33617),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__6765 (
            .O(N__33614),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__6764 (
            .O(N__33609),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__6763 (
            .O(N__33606),
            .I(N__33599));
    InMux I__6762 (
            .O(N__33605),
            .I(N__33599));
    InMux I__6761 (
            .O(N__33604),
            .I(N__33596));
    LocalMux I__6760 (
            .O(N__33599),
            .I(N__33593));
    LocalMux I__6759 (
            .O(N__33596),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__6758 (
            .O(N__33593),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__6757 (
            .O(N__33588),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__6756 (
            .O(N__33585),
            .I(N__33578));
    InMux I__6755 (
            .O(N__33584),
            .I(N__33578));
    InMux I__6754 (
            .O(N__33583),
            .I(N__33575));
    LocalMux I__6753 (
            .O(N__33578),
            .I(N__33572));
    LocalMux I__6752 (
            .O(N__33575),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__6751 (
            .O(N__33572),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__6750 (
            .O(N__33567),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__6749 (
            .O(N__33564),
            .I(N__33560));
    CascadeMux I__6748 (
            .O(N__33563),
            .I(N__33557));
    InMux I__6747 (
            .O(N__33560),
            .I(N__33551));
    InMux I__6746 (
            .O(N__33557),
            .I(N__33551));
    InMux I__6745 (
            .O(N__33556),
            .I(N__33548));
    LocalMux I__6744 (
            .O(N__33551),
            .I(N__33545));
    LocalMux I__6743 (
            .O(N__33548),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__6742 (
            .O(N__33545),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__6741 (
            .O(N__33540),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__6740 (
            .O(N__33537),
            .I(N__33534));
    InMux I__6739 (
            .O(N__33534),
            .I(N__33530));
    InMux I__6738 (
            .O(N__33533),
            .I(N__33526));
    LocalMux I__6737 (
            .O(N__33530),
            .I(N__33523));
    InMux I__6736 (
            .O(N__33529),
            .I(N__33520));
    LocalMux I__6735 (
            .O(N__33526),
            .I(N__33517));
    Span4Mux_h I__6734 (
            .O(N__33523),
            .I(N__33514));
    LocalMux I__6733 (
            .O(N__33520),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__6732 (
            .O(N__33517),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__6731 (
            .O(N__33514),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__6730 (
            .O(N__33507),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__6729 (
            .O(N__33504),
            .I(N__33498));
    InMux I__6728 (
            .O(N__33503),
            .I(N__33498));
    LocalMux I__6727 (
            .O(N__33498),
            .I(N__33494));
    InMux I__6726 (
            .O(N__33497),
            .I(N__33491));
    Span4Mux_h I__6725 (
            .O(N__33494),
            .I(N__33488));
    LocalMux I__6724 (
            .O(N__33491),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__6723 (
            .O(N__33488),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__6722 (
            .O(N__33483),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__6721 (
            .O(N__33480),
            .I(N__33477));
    InMux I__6720 (
            .O(N__33477),
            .I(N__33472));
    CascadeMux I__6719 (
            .O(N__33476),
            .I(N__33469));
    InMux I__6718 (
            .O(N__33475),
            .I(N__33466));
    LocalMux I__6717 (
            .O(N__33472),
            .I(N__33463));
    InMux I__6716 (
            .O(N__33469),
            .I(N__33460));
    LocalMux I__6715 (
            .O(N__33466),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__6714 (
            .O(N__33463),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__6713 (
            .O(N__33460),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__6712 (
            .O(N__33453),
            .I(bfn_14_14_0_));
    InMux I__6711 (
            .O(N__33450),
            .I(N__33447));
    LocalMux I__6710 (
            .O(N__33447),
            .I(N__33444));
    Odrv4 I__6709 (
            .O(N__33444),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ));
    CascadeMux I__6708 (
            .O(N__33441),
            .I(N__33436));
    InMux I__6707 (
            .O(N__33440),
            .I(N__33430));
    CascadeMux I__6706 (
            .O(N__33439),
            .I(N__33427));
    InMux I__6705 (
            .O(N__33436),
            .I(N__33422));
    InMux I__6704 (
            .O(N__33435),
            .I(N__33422));
    InMux I__6703 (
            .O(N__33434),
            .I(N__33419));
    InMux I__6702 (
            .O(N__33433),
            .I(N__33416));
    LocalMux I__6701 (
            .O(N__33430),
            .I(N__33413));
    InMux I__6700 (
            .O(N__33427),
            .I(N__33410));
    LocalMux I__6699 (
            .O(N__33422),
            .I(N__33405));
    LocalMux I__6698 (
            .O(N__33419),
            .I(N__33405));
    LocalMux I__6697 (
            .O(N__33416),
            .I(N__33402));
    Span4Mux_h I__6696 (
            .O(N__33413),
            .I(N__33397));
    LocalMux I__6695 (
            .O(N__33410),
            .I(N__33397));
    Span4Mux_h I__6694 (
            .O(N__33405),
            .I(N__33394));
    Odrv4 I__6693 (
            .O(N__33402),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    Odrv4 I__6692 (
            .O(N__33397),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    Odrv4 I__6691 (
            .O(N__33394),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ));
    CascadeMux I__6690 (
            .O(N__33387),
            .I(\delay_measurement_inst.N_360_cascade_ ));
    InMux I__6689 (
            .O(N__33384),
            .I(N__33381));
    LocalMux I__6688 (
            .O(N__33381),
            .I(N__33378));
    Span4Mux_v I__6687 (
            .O(N__33378),
            .I(N__33373));
    InMux I__6686 (
            .O(N__33377),
            .I(N__33370));
    InMux I__6685 (
            .O(N__33376),
            .I(N__33367));
    Odrv4 I__6684 (
            .O(N__33373),
            .I(measured_delay_tr_9));
    LocalMux I__6683 (
            .O(N__33370),
            .I(measured_delay_tr_9));
    LocalMux I__6682 (
            .O(N__33367),
            .I(measured_delay_tr_9));
    CascadeMux I__6681 (
            .O(N__33360),
            .I(\delay_measurement_inst.N_354_cascade_ ));
    InMux I__6680 (
            .O(N__33357),
            .I(N__33353));
    InMux I__6679 (
            .O(N__33356),
            .I(N__33350));
    LocalMux I__6678 (
            .O(N__33353),
            .I(N__33347));
    LocalMux I__6677 (
            .O(N__33350),
            .I(N__33344));
    Span4Mux_h I__6676 (
            .O(N__33347),
            .I(N__33340));
    Span4Mux_v I__6675 (
            .O(N__33344),
            .I(N__33337));
    InMux I__6674 (
            .O(N__33343),
            .I(N__33334));
    Odrv4 I__6673 (
            .O(N__33340),
            .I(measured_delay_tr_10));
    Odrv4 I__6672 (
            .O(N__33337),
            .I(measured_delay_tr_10));
    LocalMux I__6671 (
            .O(N__33334),
            .I(measured_delay_tr_10));
    InMux I__6670 (
            .O(N__33327),
            .I(N__33324));
    LocalMux I__6669 (
            .O(N__33324),
            .I(N__33321));
    Span4Mux_h I__6668 (
            .O(N__33321),
            .I(N__33316));
    InMux I__6667 (
            .O(N__33320),
            .I(N__33313));
    InMux I__6666 (
            .O(N__33319),
            .I(N__33310));
    Odrv4 I__6665 (
            .O(N__33316),
            .I(measured_delay_tr_11));
    LocalMux I__6664 (
            .O(N__33313),
            .I(measured_delay_tr_11));
    LocalMux I__6663 (
            .O(N__33310),
            .I(measured_delay_tr_11));
    InMux I__6662 (
            .O(N__33303),
            .I(N__33299));
    InMux I__6661 (
            .O(N__33302),
            .I(N__33296));
    LocalMux I__6660 (
            .O(N__33299),
            .I(N__33293));
    LocalMux I__6659 (
            .O(N__33296),
            .I(N__33290));
    Span4Mux_h I__6658 (
            .O(N__33293),
            .I(N__33286));
    Span4Mux_h I__6657 (
            .O(N__33290),
            .I(N__33283));
    InMux I__6656 (
            .O(N__33289),
            .I(N__33280));
    Odrv4 I__6655 (
            .O(N__33286),
            .I(measured_delay_tr_12));
    Odrv4 I__6654 (
            .O(N__33283),
            .I(measured_delay_tr_12));
    LocalMux I__6653 (
            .O(N__33280),
            .I(measured_delay_tr_12));
    InMux I__6652 (
            .O(N__33273),
            .I(N__33261));
    InMux I__6651 (
            .O(N__33272),
            .I(N__33261));
    InMux I__6650 (
            .O(N__33271),
            .I(N__33261));
    InMux I__6649 (
            .O(N__33270),
            .I(N__33261));
    LocalMux I__6648 (
            .O(N__33261),
            .I(\delay_measurement_inst.N_354 ));
    InMux I__6647 (
            .O(N__33258),
            .I(N__33254));
    InMux I__6646 (
            .O(N__33257),
            .I(N__33251));
    LocalMux I__6645 (
            .O(N__33254),
            .I(N__33245));
    LocalMux I__6644 (
            .O(N__33251),
            .I(N__33245));
    CascadeMux I__6643 (
            .O(N__33250),
            .I(N__33242));
    Span4Mux_h I__6642 (
            .O(N__33245),
            .I(N__33239));
    InMux I__6641 (
            .O(N__33242),
            .I(N__33236));
    Odrv4 I__6640 (
            .O(N__33239),
            .I(measured_delay_tr_13));
    LocalMux I__6639 (
            .O(N__33236),
            .I(measured_delay_tr_13));
    InMux I__6638 (
            .O(N__33231),
            .I(N__33228));
    LocalMux I__6637 (
            .O(N__33228),
            .I(N__33224));
    InMux I__6636 (
            .O(N__33227),
            .I(N__33221));
    Span12Mux_v I__6635 (
            .O(N__33224),
            .I(N__33218));
    LocalMux I__6634 (
            .O(N__33221),
            .I(N__33215));
    Span12Mux_h I__6633 (
            .O(N__33218),
            .I(N__33212));
    Span4Mux_s2_h I__6632 (
            .O(N__33215),
            .I(N__33209));
    Odrv12 I__6631 (
            .O(N__33212),
            .I(pwm_duty_input_1));
    Odrv4 I__6630 (
            .O(N__33209),
            .I(pwm_duty_input_1));
    InMux I__6629 (
            .O(N__33204),
            .I(N__33201));
    LocalMux I__6628 (
            .O(N__33201),
            .I(N__33197));
    InMux I__6627 (
            .O(N__33200),
            .I(N__33194));
    Span12Mux_v I__6626 (
            .O(N__33197),
            .I(N__33191));
    LocalMux I__6625 (
            .O(N__33194),
            .I(N__33188));
    Span12Mux_h I__6624 (
            .O(N__33191),
            .I(N__33185));
    Span4Mux_v I__6623 (
            .O(N__33188),
            .I(N__33182));
    Odrv12 I__6622 (
            .O(N__33185),
            .I(pwm_duty_input_0));
    Odrv4 I__6621 (
            .O(N__33182),
            .I(pwm_duty_input_0));
    InMux I__6620 (
            .O(N__33177),
            .I(N__33174));
    LocalMux I__6619 (
            .O(N__33174),
            .I(N__33171));
    Span4Mux_v I__6618 (
            .O(N__33171),
            .I(N__33167));
    InMux I__6617 (
            .O(N__33170),
            .I(N__33164));
    Span4Mux_h I__6616 (
            .O(N__33167),
            .I(N__33161));
    LocalMux I__6615 (
            .O(N__33164),
            .I(N__33158));
    Sp12to4 I__6614 (
            .O(N__33161),
            .I(N__33155));
    Span4Mux_v I__6613 (
            .O(N__33158),
            .I(N__33152));
    Odrv12 I__6612 (
            .O(N__33155),
            .I(pwm_duty_input_2));
    Odrv4 I__6611 (
            .O(N__33152),
            .I(pwm_duty_input_2));
    InMux I__6610 (
            .O(N__33147),
            .I(N__33144));
    LocalMux I__6609 (
            .O(N__33144),
            .I(N__33141));
    Span12Mux_s8_h I__6608 (
            .O(N__33141),
            .I(N__33138));
    Odrv12 I__6607 (
            .O(N__33138),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    CascadeMux I__6606 (
            .O(N__33135),
            .I(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ));
    CascadeMux I__6605 (
            .O(N__33132),
            .I(N__33128));
    CascadeMux I__6604 (
            .O(N__33131),
            .I(N__33124));
    InMux I__6603 (
            .O(N__33128),
            .I(N__33121));
    InMux I__6602 (
            .O(N__33127),
            .I(N__33118));
    InMux I__6601 (
            .O(N__33124),
            .I(N__33115));
    LocalMux I__6600 (
            .O(N__33121),
            .I(N__33110));
    LocalMux I__6599 (
            .O(N__33118),
            .I(N__33110));
    LocalMux I__6598 (
            .O(N__33115),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    Odrv4 I__6597 (
            .O(N__33110),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ));
    CascadeMux I__6596 (
            .O(N__33105),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ));
    InMux I__6595 (
            .O(N__33102),
            .I(N__33098));
    InMux I__6594 (
            .O(N__33101),
            .I(N__33095));
    LocalMux I__6593 (
            .O(N__33098),
            .I(N__33092));
    LocalMux I__6592 (
            .O(N__33095),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    Odrv4 I__6591 (
            .O(N__33092),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ));
    InMux I__6590 (
            .O(N__33087),
            .I(N__33084));
    LocalMux I__6589 (
            .O(N__33084),
            .I(N__33081));
    Span4Mux_v I__6588 (
            .O(N__33081),
            .I(N__33078));
    Odrv4 I__6587 (
            .O(N__33078),
            .I(delay_tr_input_c));
    InMux I__6586 (
            .O(N__33075),
            .I(N__33072));
    LocalMux I__6585 (
            .O(N__33072),
            .I(delay_tr_d1));
    InMux I__6584 (
            .O(N__33069),
            .I(N__33063));
    InMux I__6583 (
            .O(N__33068),
            .I(N__33063));
    LocalMux I__6582 (
            .O(N__33063),
            .I(N__33058));
    InMux I__6581 (
            .O(N__33062),
            .I(N__33055));
    InMux I__6580 (
            .O(N__33061),
            .I(N__33052));
    Span4Mux_v I__6579 (
            .O(N__33058),
            .I(N__33047));
    LocalMux I__6578 (
            .O(N__33055),
            .I(N__33047));
    LocalMux I__6577 (
            .O(N__33052),
            .I(delay_tr_d2));
    Odrv4 I__6576 (
            .O(N__33047),
            .I(delay_tr_d2));
    InMux I__6575 (
            .O(N__33042),
            .I(N__33039));
    LocalMux I__6574 (
            .O(N__33039),
            .I(N__33036));
    Span4Mux_h I__6573 (
            .O(N__33036),
            .I(N__33033));
    Span4Mux_h I__6572 (
            .O(N__33033),
            .I(N__33030));
    Sp12to4 I__6571 (
            .O(N__33030),
            .I(N__33027));
    Odrv12 I__6570 (
            .O(N__33027),
            .I(il_min_comp1_c));
    CascadeMux I__6569 (
            .O(N__33024),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    IoInMux I__6568 (
            .O(N__33021),
            .I(N__33018));
    LocalMux I__6567 (
            .O(N__33018),
            .I(N__33015));
    Span4Mux_s1_v I__6566 (
            .O(N__33015),
            .I(N__33012));
    Span4Mux_v I__6565 (
            .O(N__33012),
            .I(N__33009));
    Span4Mux_v I__6564 (
            .O(N__33009),
            .I(N__33004));
    InMux I__6563 (
            .O(N__33008),
            .I(N__32999));
    InMux I__6562 (
            .O(N__33007),
            .I(N__32999));
    Odrv4 I__6561 (
            .O(N__33004),
            .I(s1_phy_c));
    LocalMux I__6560 (
            .O(N__32999),
            .I(s1_phy_c));
    InMux I__6559 (
            .O(N__32994),
            .I(N__32990));
    InMux I__6558 (
            .O(N__32993),
            .I(N__32987));
    LocalMux I__6557 (
            .O(N__32990),
            .I(N__32982));
    LocalMux I__6556 (
            .O(N__32987),
            .I(N__32982));
    Span4Mux_h I__6555 (
            .O(N__32982),
            .I(N__32979));
    Span4Mux_v I__6554 (
            .O(N__32979),
            .I(N__32975));
    InMux I__6553 (
            .O(N__32978),
            .I(N__32972));
    Odrv4 I__6552 (
            .O(N__32975),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    LocalMux I__6551 (
            .O(N__32972),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__6550 (
            .O(N__32967),
            .I(N__32946));
    CEMux I__6549 (
            .O(N__32966),
            .I(N__32946));
    CEMux I__6548 (
            .O(N__32965),
            .I(N__32946));
    CEMux I__6547 (
            .O(N__32964),
            .I(N__32946));
    CEMux I__6546 (
            .O(N__32963),
            .I(N__32946));
    CEMux I__6545 (
            .O(N__32962),
            .I(N__32946));
    CEMux I__6544 (
            .O(N__32961),
            .I(N__32946));
    GlobalMux I__6543 (
            .O(N__32946),
            .I(N__32943));
    gio2CtrlBuf I__6542 (
            .O(N__32943),
            .I(\current_shift_inst.timer_s1.N_185_i_g ));
    InMux I__6541 (
            .O(N__32940),
            .I(N__32936));
    InMux I__6540 (
            .O(N__32939),
            .I(N__32933));
    LocalMux I__6539 (
            .O(N__32936),
            .I(N__32927));
    LocalMux I__6538 (
            .O(N__32933),
            .I(N__32927));
    InMux I__6537 (
            .O(N__32932),
            .I(N__32924));
    Span4Mux_v I__6536 (
            .O(N__32927),
            .I(N__32918));
    LocalMux I__6535 (
            .O(N__32924),
            .I(N__32918));
    InMux I__6534 (
            .O(N__32923),
            .I(N__32915));
    Odrv4 I__6533 (
            .O(N__32918),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__6532 (
            .O(N__32915),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__6531 (
            .O(N__32910),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__6530 (
            .O(N__32907),
            .I(N__32903));
    InMux I__6529 (
            .O(N__32906),
            .I(N__32900));
    LocalMux I__6528 (
            .O(N__32903),
            .I(N__32896));
    LocalMux I__6527 (
            .O(N__32900),
            .I(N__32893));
    InMux I__6526 (
            .O(N__32899),
            .I(N__32890));
    Span4Mux_h I__6525 (
            .O(N__32896),
            .I(N__32886));
    Span4Mux_v I__6524 (
            .O(N__32893),
            .I(N__32881));
    LocalMux I__6523 (
            .O(N__32890),
            .I(N__32881));
    InMux I__6522 (
            .O(N__32889),
            .I(N__32878));
    Odrv4 I__6521 (
            .O(N__32886),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__6520 (
            .O(N__32881),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__6519 (
            .O(N__32878),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__6518 (
            .O(N__32871),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__6517 (
            .O(N__32868),
            .I(N__32864));
    InMux I__6516 (
            .O(N__32867),
            .I(N__32860));
    LocalMux I__6515 (
            .O(N__32864),
            .I(N__32857));
    InMux I__6514 (
            .O(N__32863),
            .I(N__32853));
    LocalMux I__6513 (
            .O(N__32860),
            .I(N__32850));
    Sp12to4 I__6512 (
            .O(N__32857),
            .I(N__32847));
    InMux I__6511 (
            .O(N__32856),
            .I(N__32844));
    LocalMux I__6510 (
            .O(N__32853),
            .I(N__32841));
    Span4Mux_h I__6509 (
            .O(N__32850),
            .I(N__32838));
    Span12Mux_v I__6508 (
            .O(N__32847),
            .I(N__32831));
    LocalMux I__6507 (
            .O(N__32844),
            .I(N__32831));
    Span12Mux_v I__6506 (
            .O(N__32841),
            .I(N__32831));
    Odrv4 I__6505 (
            .O(N__32838),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__6504 (
            .O(N__32831),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__6503 (
            .O(N__32826),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__6502 (
            .O(N__32823),
            .I(N__32820));
    InMux I__6501 (
            .O(N__32820),
            .I(N__32813));
    InMux I__6500 (
            .O(N__32819),
            .I(N__32813));
    InMux I__6499 (
            .O(N__32818),
            .I(N__32810));
    LocalMux I__6498 (
            .O(N__32813),
            .I(N__32807));
    LocalMux I__6497 (
            .O(N__32810),
            .I(N__32804));
    Span4Mux_v I__6496 (
            .O(N__32807),
            .I(N__32800));
    Span4Mux_h I__6495 (
            .O(N__32804),
            .I(N__32797));
    InMux I__6494 (
            .O(N__32803),
            .I(N__32794));
    Odrv4 I__6493 (
            .O(N__32800),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__6492 (
            .O(N__32797),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__6491 (
            .O(N__32794),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__6490 (
            .O(N__32787),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__6489 (
            .O(N__32784),
            .I(N__32780));
    InMux I__6488 (
            .O(N__32783),
            .I(N__32772));
    InMux I__6487 (
            .O(N__32780),
            .I(N__32772));
    InMux I__6486 (
            .O(N__32779),
            .I(N__32772));
    LocalMux I__6485 (
            .O(N__32772),
            .I(N__32768));
    InMux I__6484 (
            .O(N__32771),
            .I(N__32765));
    Odrv4 I__6483 (
            .O(N__32768),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__6482 (
            .O(N__32765),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__6481 (
            .O(N__32760),
            .I(bfn_13_18_0_));
    InMux I__6480 (
            .O(N__32757),
            .I(N__32753));
    CascadeMux I__6479 (
            .O(N__32756),
            .I(N__32750));
    LocalMux I__6478 (
            .O(N__32753),
            .I(N__32746));
    InMux I__6477 (
            .O(N__32750),
            .I(N__32741));
    InMux I__6476 (
            .O(N__32749),
            .I(N__32741));
    Span12Mux_v I__6475 (
            .O(N__32746),
            .I(N__32735));
    LocalMux I__6474 (
            .O(N__32741),
            .I(N__32735));
    InMux I__6473 (
            .O(N__32740),
            .I(N__32732));
    Odrv12 I__6472 (
            .O(N__32735),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__6471 (
            .O(N__32732),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__6470 (
            .O(N__32727),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__6469 (
            .O(N__32724),
            .I(N__32720));
    CascadeMux I__6468 (
            .O(N__32723),
            .I(N__32717));
    LocalMux I__6467 (
            .O(N__32720),
            .I(N__32713));
    InMux I__6466 (
            .O(N__32717),
            .I(N__32708));
    InMux I__6465 (
            .O(N__32716),
            .I(N__32708));
    Span4Mux_h I__6464 (
            .O(N__32713),
            .I(N__32704));
    LocalMux I__6463 (
            .O(N__32708),
            .I(N__32701));
    InMux I__6462 (
            .O(N__32707),
            .I(N__32698));
    Odrv4 I__6461 (
            .O(N__32704),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__6460 (
            .O(N__32701),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__6459 (
            .O(N__32698),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__6458 (
            .O(N__32691),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__6457 (
            .O(N__32688),
            .I(N__32684));
    InMux I__6456 (
            .O(N__32687),
            .I(N__32681));
    LocalMux I__6455 (
            .O(N__32684),
            .I(N__32676));
    LocalMux I__6454 (
            .O(N__32681),
            .I(N__32673));
    InMux I__6453 (
            .O(N__32680),
            .I(N__32670));
    InMux I__6452 (
            .O(N__32679),
            .I(N__32667));
    Span4Mux_h I__6451 (
            .O(N__32676),
            .I(N__32664));
    Span4Mux_v I__6450 (
            .O(N__32673),
            .I(N__32657));
    LocalMux I__6449 (
            .O(N__32670),
            .I(N__32657));
    LocalMux I__6448 (
            .O(N__32667),
            .I(N__32657));
    Odrv4 I__6447 (
            .O(N__32664),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__6446 (
            .O(N__32657),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__6445 (
            .O(N__32652),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__6444 (
            .O(N__32649),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__6443 (
            .O(N__32646),
            .I(N__32641));
    InMux I__6442 (
            .O(N__32645),
            .I(N__32638));
    InMux I__6441 (
            .O(N__32644),
            .I(N__32635));
    LocalMux I__6440 (
            .O(N__32641),
            .I(N__32630));
    LocalMux I__6439 (
            .O(N__32638),
            .I(N__32630));
    LocalMux I__6438 (
            .O(N__32635),
            .I(N__32627));
    Span4Mux_v I__6437 (
            .O(N__32630),
            .I(N__32623));
    Span4Mux_h I__6436 (
            .O(N__32627),
            .I(N__32620));
    InMux I__6435 (
            .O(N__32626),
            .I(N__32617));
    Odrv4 I__6434 (
            .O(N__32623),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__6433 (
            .O(N__32620),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__6432 (
            .O(N__32617),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__6431 (
            .O(N__32610),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__6430 (
            .O(N__32607),
            .I(N__32602));
    InMux I__6429 (
            .O(N__32606),
            .I(N__32599));
    InMux I__6428 (
            .O(N__32605),
            .I(N__32596));
    LocalMux I__6427 (
            .O(N__32602),
            .I(N__32591));
    LocalMux I__6426 (
            .O(N__32599),
            .I(N__32591));
    LocalMux I__6425 (
            .O(N__32596),
            .I(N__32588));
    Span4Mux_v I__6424 (
            .O(N__32591),
            .I(N__32584));
    Span4Mux_h I__6423 (
            .O(N__32588),
            .I(N__32581));
    InMux I__6422 (
            .O(N__32587),
            .I(N__32578));
    Odrv4 I__6421 (
            .O(N__32584),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__6420 (
            .O(N__32581),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__6419 (
            .O(N__32578),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__6418 (
            .O(N__32571),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__6417 (
            .O(N__32568),
            .I(N__32562));
    InMux I__6416 (
            .O(N__32567),
            .I(N__32559));
    InMux I__6415 (
            .O(N__32566),
            .I(N__32556));
    InMux I__6414 (
            .O(N__32565),
            .I(N__32553));
    LocalMux I__6413 (
            .O(N__32562),
            .I(N__32550));
    LocalMux I__6412 (
            .O(N__32559),
            .I(N__32545));
    LocalMux I__6411 (
            .O(N__32556),
            .I(N__32545));
    LocalMux I__6410 (
            .O(N__32553),
            .I(N__32542));
    Span4Mux_h I__6409 (
            .O(N__32550),
            .I(N__32539));
    Span12Mux_v I__6408 (
            .O(N__32545),
            .I(N__32534));
    Span12Mux_v I__6407 (
            .O(N__32542),
            .I(N__32534));
    Odrv4 I__6406 (
            .O(N__32539),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv12 I__6405 (
            .O(N__32534),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__6404 (
            .O(N__32529),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__6403 (
            .O(N__32526),
            .I(N__32523));
    LocalMux I__6402 (
            .O(N__32523),
            .I(N__32518));
    InMux I__6401 (
            .O(N__32522),
            .I(N__32515));
    InMux I__6400 (
            .O(N__32521),
            .I(N__32512));
    Span4Mux_h I__6399 (
            .O(N__32518),
            .I(N__32506));
    LocalMux I__6398 (
            .O(N__32515),
            .I(N__32506));
    LocalMux I__6397 (
            .O(N__32512),
            .I(N__32503));
    InMux I__6396 (
            .O(N__32511),
            .I(N__32500));
    Span4Mux_v I__6395 (
            .O(N__32506),
            .I(N__32495));
    Span4Mux_h I__6394 (
            .O(N__32503),
            .I(N__32495));
    LocalMux I__6393 (
            .O(N__32500),
            .I(N__32492));
    Odrv4 I__6392 (
            .O(N__32495),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv12 I__6391 (
            .O(N__32492),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__6390 (
            .O(N__32487),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__6389 (
            .O(N__32484),
            .I(N__32481));
    LocalMux I__6388 (
            .O(N__32481),
            .I(N__32477));
    CascadeMux I__6387 (
            .O(N__32480),
            .I(N__32474));
    Sp12to4 I__6386 (
            .O(N__32477),
            .I(N__32470));
    InMux I__6385 (
            .O(N__32474),
            .I(N__32465));
    InMux I__6384 (
            .O(N__32473),
            .I(N__32465));
    Span12Mux_v I__6383 (
            .O(N__32470),
            .I(N__32459));
    LocalMux I__6382 (
            .O(N__32465),
            .I(N__32459));
    InMux I__6381 (
            .O(N__32464),
            .I(N__32456));
    Odrv12 I__6380 (
            .O(N__32459),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__6379 (
            .O(N__32456),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__6378 (
            .O(N__32451),
            .I(bfn_13_17_0_));
    InMux I__6377 (
            .O(N__32448),
            .I(N__32443));
    InMux I__6376 (
            .O(N__32447),
            .I(N__32440));
    InMux I__6375 (
            .O(N__32446),
            .I(N__32437));
    LocalMux I__6374 (
            .O(N__32443),
            .I(N__32432));
    LocalMux I__6373 (
            .O(N__32440),
            .I(N__32432));
    LocalMux I__6372 (
            .O(N__32437),
            .I(N__32429));
    Span4Mux_v I__6371 (
            .O(N__32432),
            .I(N__32423));
    Span4Mux_v I__6370 (
            .O(N__32429),
            .I(N__32423));
    InMux I__6369 (
            .O(N__32428),
            .I(N__32420));
    Odrv4 I__6368 (
            .O(N__32423),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__6367 (
            .O(N__32420),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__6366 (
            .O(N__32415),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__6365 (
            .O(N__32412),
            .I(N__32408));
    InMux I__6364 (
            .O(N__32411),
            .I(N__32405));
    LocalMux I__6363 (
            .O(N__32408),
            .I(N__32401));
    LocalMux I__6362 (
            .O(N__32405),
            .I(N__32398));
    InMux I__6361 (
            .O(N__32404),
            .I(N__32395));
    Span4Mux_h I__6360 (
            .O(N__32401),
            .I(N__32391));
    Span4Mux_v I__6359 (
            .O(N__32398),
            .I(N__32386));
    LocalMux I__6358 (
            .O(N__32395),
            .I(N__32386));
    InMux I__6357 (
            .O(N__32394),
            .I(N__32383));
    Odrv4 I__6356 (
            .O(N__32391),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__6355 (
            .O(N__32386),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__6354 (
            .O(N__32383),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__6353 (
            .O(N__32376),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__6352 (
            .O(N__32373),
            .I(N__32370));
    LocalMux I__6351 (
            .O(N__32370),
            .I(N__32366));
    InMux I__6350 (
            .O(N__32369),
            .I(N__32363));
    Span4Mux_h I__6349 (
            .O(N__32366),
            .I(N__32358));
    LocalMux I__6348 (
            .O(N__32363),
            .I(N__32358));
    Span4Mux_v I__6347 (
            .O(N__32358),
            .I(N__32353));
    InMux I__6346 (
            .O(N__32357),
            .I(N__32350));
    InMux I__6345 (
            .O(N__32356),
            .I(N__32347));
    Odrv4 I__6344 (
            .O(N__32353),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__6343 (
            .O(N__32350),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__6342 (
            .O(N__32347),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__6341 (
            .O(N__32340),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__6340 (
            .O(N__32337),
            .I(N__32333));
    CascadeMux I__6339 (
            .O(N__32336),
            .I(N__32329));
    InMux I__6338 (
            .O(N__32333),
            .I(N__32326));
    InMux I__6337 (
            .O(N__32332),
            .I(N__32323));
    InMux I__6336 (
            .O(N__32329),
            .I(N__32320));
    LocalMux I__6335 (
            .O(N__32326),
            .I(N__32317));
    LocalMux I__6334 (
            .O(N__32323),
            .I(N__32314));
    LocalMux I__6333 (
            .O(N__32320),
            .I(N__32308));
    Span4Mux_h I__6332 (
            .O(N__32317),
            .I(N__32308));
    Span4Mux_h I__6331 (
            .O(N__32314),
            .I(N__32305));
    InMux I__6330 (
            .O(N__32313),
            .I(N__32302));
    Odrv4 I__6329 (
            .O(N__32308),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__6328 (
            .O(N__32305),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__6327 (
            .O(N__32302),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__6326 (
            .O(N__32295),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__6325 (
            .O(N__32292),
            .I(N__32288));
    InMux I__6324 (
            .O(N__32291),
            .I(N__32284));
    LocalMux I__6323 (
            .O(N__32288),
            .I(N__32281));
    InMux I__6322 (
            .O(N__32287),
            .I(N__32278));
    LocalMux I__6321 (
            .O(N__32284),
            .I(N__32275));
    Span4Mux_h I__6320 (
            .O(N__32281),
            .I(N__32272));
    LocalMux I__6319 (
            .O(N__32278),
            .I(N__32269));
    Span4Mux_v I__6318 (
            .O(N__32275),
            .I(N__32265));
    Span4Mux_h I__6317 (
            .O(N__32272),
            .I(N__32260));
    Span4Mux_h I__6316 (
            .O(N__32269),
            .I(N__32260));
    InMux I__6315 (
            .O(N__32268),
            .I(N__32257));
    Odrv4 I__6314 (
            .O(N__32265),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__6313 (
            .O(N__32260),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__6312 (
            .O(N__32257),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__6311 (
            .O(N__32250),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__6310 (
            .O(N__32247),
            .I(N__32244));
    LocalMux I__6309 (
            .O(N__32244),
            .I(N__32240));
    InMux I__6308 (
            .O(N__32243),
            .I(N__32237));
    Span4Mux_v I__6307 (
            .O(N__32240),
            .I(N__32231));
    LocalMux I__6306 (
            .O(N__32237),
            .I(N__32231));
    InMux I__6305 (
            .O(N__32236),
            .I(N__32228));
    Span4Mux_v I__6304 (
            .O(N__32231),
            .I(N__32224));
    LocalMux I__6303 (
            .O(N__32228),
            .I(N__32221));
    InMux I__6302 (
            .O(N__32227),
            .I(N__32218));
    Odrv4 I__6301 (
            .O(N__32224),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__6300 (
            .O(N__32221),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__6299 (
            .O(N__32218),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__6298 (
            .O(N__32211),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__6297 (
            .O(N__32208),
            .I(N__32205));
    InMux I__6296 (
            .O(N__32205),
            .I(N__32201));
    InMux I__6295 (
            .O(N__32204),
            .I(N__32198));
    LocalMux I__6294 (
            .O(N__32201),
            .I(N__32194));
    LocalMux I__6293 (
            .O(N__32198),
            .I(N__32191));
    InMux I__6292 (
            .O(N__32197),
            .I(N__32188));
    Span4Mux_v I__6291 (
            .O(N__32194),
            .I(N__32180));
    Span4Mux_v I__6290 (
            .O(N__32191),
            .I(N__32180));
    LocalMux I__6289 (
            .O(N__32188),
            .I(N__32180));
    InMux I__6288 (
            .O(N__32187),
            .I(N__32177));
    Odrv4 I__6287 (
            .O(N__32180),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__6286 (
            .O(N__32177),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__6285 (
            .O(N__32172),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__6284 (
            .O(N__32169),
            .I(N__32164));
    InMux I__6283 (
            .O(N__32168),
            .I(N__32161));
    InMux I__6282 (
            .O(N__32167),
            .I(N__32158));
    LocalMux I__6281 (
            .O(N__32164),
            .I(N__32155));
    LocalMux I__6280 (
            .O(N__32161),
            .I(N__32152));
    LocalMux I__6279 (
            .O(N__32158),
            .I(N__32149));
    Span4Mux_v I__6278 (
            .O(N__32155),
            .I(N__32145));
    Span4Mux_v I__6277 (
            .O(N__32152),
            .I(N__32140));
    Span4Mux_h I__6276 (
            .O(N__32149),
            .I(N__32140));
    InMux I__6275 (
            .O(N__32148),
            .I(N__32137));
    Odrv4 I__6274 (
            .O(N__32145),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__6273 (
            .O(N__32140),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__6272 (
            .O(N__32137),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__6271 (
            .O(N__32130),
            .I(bfn_13_16_0_));
    CascadeMux I__6270 (
            .O(N__32127),
            .I(N__32123));
    InMux I__6269 (
            .O(N__32126),
            .I(N__32120));
    InMux I__6268 (
            .O(N__32123),
            .I(N__32116));
    LocalMux I__6267 (
            .O(N__32120),
            .I(N__32113));
    InMux I__6266 (
            .O(N__32119),
            .I(N__32110));
    LocalMux I__6265 (
            .O(N__32116),
            .I(N__32105));
    Span4Mux_v I__6264 (
            .O(N__32113),
            .I(N__32105));
    LocalMux I__6263 (
            .O(N__32110),
            .I(N__32102));
    Span4Mux_v I__6262 (
            .O(N__32105),
            .I(N__32096));
    Span4Mux_v I__6261 (
            .O(N__32102),
            .I(N__32096));
    InMux I__6260 (
            .O(N__32101),
            .I(N__32093));
    Odrv4 I__6259 (
            .O(N__32096),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__6258 (
            .O(N__32093),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__6257 (
            .O(N__32088),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__6256 (
            .O(N__32085),
            .I(N__32081));
    InMux I__6255 (
            .O(N__32084),
            .I(N__32077));
    LocalMux I__6254 (
            .O(N__32081),
            .I(N__32074));
    InMux I__6253 (
            .O(N__32080),
            .I(N__32071));
    LocalMux I__6252 (
            .O(N__32077),
            .I(N__32068));
    Span4Mux_v I__6251 (
            .O(N__32074),
            .I(N__32062));
    LocalMux I__6250 (
            .O(N__32071),
            .I(N__32062));
    Span4Mux_h I__6249 (
            .O(N__32068),
            .I(N__32059));
    InMux I__6248 (
            .O(N__32067),
            .I(N__32056));
    Odrv4 I__6247 (
            .O(N__32062),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__6246 (
            .O(N__32059),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__6245 (
            .O(N__32056),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__6244 (
            .O(N__32049),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__6243 (
            .O(N__32046),
            .I(N__32042));
    InMux I__6242 (
            .O(N__32045),
            .I(N__32038));
    LocalMux I__6241 (
            .O(N__32042),
            .I(N__32035));
    InMux I__6240 (
            .O(N__32041),
            .I(N__32032));
    LocalMux I__6239 (
            .O(N__32038),
            .I(N__32029));
    Span4Mux_h I__6238 (
            .O(N__32035),
            .I(N__32026));
    LocalMux I__6237 (
            .O(N__32032),
            .I(N__32023));
    Span4Mux_h I__6236 (
            .O(N__32029),
            .I(N__32019));
    Span4Mux_v I__6235 (
            .O(N__32026),
            .I(N__32014));
    Span4Mux_h I__6234 (
            .O(N__32023),
            .I(N__32014));
    InMux I__6233 (
            .O(N__32022),
            .I(N__32011));
    Odrv4 I__6232 (
            .O(N__32019),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__6231 (
            .O(N__32014),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__6230 (
            .O(N__32011),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__6229 (
            .O(N__32004),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__6228 (
            .O(N__32001),
            .I(N__31993));
    InMux I__6227 (
            .O(N__32000),
            .I(N__31988));
    InMux I__6226 (
            .O(N__31999),
            .I(N__31988));
    InMux I__6225 (
            .O(N__31998),
            .I(N__31983));
    InMux I__6224 (
            .O(N__31997),
            .I(N__31983));
    InMux I__6223 (
            .O(N__31996),
            .I(N__31980));
    LocalMux I__6222 (
            .O(N__31993),
            .I(N__31972));
    LocalMux I__6221 (
            .O(N__31988),
            .I(N__31972));
    LocalMux I__6220 (
            .O(N__31983),
            .I(N__31972));
    LocalMux I__6219 (
            .O(N__31980),
            .I(N__31968));
    InMux I__6218 (
            .O(N__31979),
            .I(N__31963));
    Span4Mux_v I__6217 (
            .O(N__31972),
            .I(N__31960));
    InMux I__6216 (
            .O(N__31971),
            .I(N__31957));
    Span4Mux_h I__6215 (
            .O(N__31968),
            .I(N__31954));
    InMux I__6214 (
            .O(N__31967),
            .I(N__31949));
    InMux I__6213 (
            .O(N__31966),
            .I(N__31949));
    LocalMux I__6212 (
            .O(N__31963),
            .I(measured_delay_tr_15));
    Odrv4 I__6211 (
            .O(N__31960),
            .I(measured_delay_tr_15));
    LocalMux I__6210 (
            .O(N__31957),
            .I(measured_delay_tr_15));
    Odrv4 I__6209 (
            .O(N__31954),
            .I(measured_delay_tr_15));
    LocalMux I__6208 (
            .O(N__31949),
            .I(measured_delay_tr_15));
    InMux I__6207 (
            .O(N__31938),
            .I(N__31933));
    InMux I__6206 (
            .O(N__31937),
            .I(N__31930));
    InMux I__6205 (
            .O(N__31936),
            .I(N__31927));
    LocalMux I__6204 (
            .O(N__31933),
            .I(N__31924));
    LocalMux I__6203 (
            .O(N__31930),
            .I(N__31919));
    LocalMux I__6202 (
            .O(N__31927),
            .I(N__31919));
    Span4Mux_h I__6201 (
            .O(N__31924),
            .I(N__31914));
    Span4Mux_h I__6200 (
            .O(N__31919),
            .I(N__31911));
    InMux I__6199 (
            .O(N__31918),
            .I(N__31908));
    InMux I__6198 (
            .O(N__31917),
            .I(N__31905));
    Odrv4 I__6197 (
            .O(N__31914),
            .I(measured_delay_tr_14));
    Odrv4 I__6196 (
            .O(N__31911),
            .I(measured_delay_tr_14));
    LocalMux I__6195 (
            .O(N__31908),
            .I(measured_delay_tr_14));
    LocalMux I__6194 (
            .O(N__31905),
            .I(measured_delay_tr_14));
    CascadeMux I__6193 (
            .O(N__31896),
            .I(N__31892));
    CascadeMux I__6192 (
            .O(N__31895),
            .I(N__31887));
    InMux I__6191 (
            .O(N__31892),
            .I(N__31870));
    InMux I__6190 (
            .O(N__31891),
            .I(N__31870));
    InMux I__6189 (
            .O(N__31890),
            .I(N__31863));
    InMux I__6188 (
            .O(N__31887),
            .I(N__31863));
    InMux I__6187 (
            .O(N__31886),
            .I(N__31863));
    InMux I__6186 (
            .O(N__31885),
            .I(N__31856));
    InMux I__6185 (
            .O(N__31884),
            .I(N__31856));
    InMux I__6184 (
            .O(N__31883),
            .I(N__31856));
    InMux I__6183 (
            .O(N__31882),
            .I(N__31847));
    InMux I__6182 (
            .O(N__31881),
            .I(N__31847));
    InMux I__6181 (
            .O(N__31880),
            .I(N__31847));
    InMux I__6180 (
            .O(N__31879),
            .I(N__31847));
    InMux I__6179 (
            .O(N__31878),
            .I(N__31838));
    InMux I__6178 (
            .O(N__31877),
            .I(N__31838));
    InMux I__6177 (
            .O(N__31876),
            .I(N__31838));
    InMux I__6176 (
            .O(N__31875),
            .I(N__31838));
    LocalMux I__6175 (
            .O(N__31870),
            .I(N__31833));
    LocalMux I__6174 (
            .O(N__31863),
            .I(N__31833));
    LocalMux I__6173 (
            .O(N__31856),
            .I(N__31830));
    LocalMux I__6172 (
            .O(N__31847),
            .I(N__31827));
    LocalMux I__6171 (
            .O(N__31838),
            .I(N__31824));
    Span4Mux_h I__6170 (
            .O(N__31833),
            .I(N__31821));
    Span4Mux_h I__6169 (
            .O(N__31830),
            .I(N__31814));
    Span4Mux_v I__6168 (
            .O(N__31827),
            .I(N__31814));
    Span4Mux_v I__6167 (
            .O(N__31824),
            .I(N__31814));
    Odrv4 I__6166 (
            .O(N__31821),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    Odrv4 I__6165 (
            .O(N__31814),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ));
    CascadeMux I__6164 (
            .O(N__31809),
            .I(N__31806));
    InMux I__6163 (
            .O(N__31806),
            .I(N__31803));
    LocalMux I__6162 (
            .O(N__31803),
            .I(\delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14 ));
    InMux I__6161 (
            .O(N__31800),
            .I(N__31797));
    LocalMux I__6160 (
            .O(N__31797),
            .I(N__31794));
    Span4Mux_v I__6159 (
            .O(N__31794),
            .I(N__31789));
    InMux I__6158 (
            .O(N__31793),
            .I(N__31786));
    InMux I__6157 (
            .O(N__31792),
            .I(N__31783));
    Span4Mux_h I__6156 (
            .O(N__31789),
            .I(N__31780));
    LocalMux I__6155 (
            .O(N__31786),
            .I(N__31777));
    LocalMux I__6154 (
            .O(N__31783),
            .I(il_min_comp2_D2));
    Odrv4 I__6153 (
            .O(N__31780),
            .I(il_min_comp2_D2));
    Odrv12 I__6152 (
            .O(N__31777),
            .I(il_min_comp2_D2));
    InMux I__6151 (
            .O(N__31770),
            .I(N__31767));
    LocalMux I__6150 (
            .O(N__31767),
            .I(N__31764));
    Span4Mux_h I__6149 (
            .O(N__31764),
            .I(N__31761));
    Span4Mux_v I__6148 (
            .O(N__31761),
            .I(N__31756));
    InMux I__6147 (
            .O(N__31760),
            .I(N__31753));
    InMux I__6146 (
            .O(N__31759),
            .I(N__31750));
    Odrv4 I__6145 (
            .O(N__31756),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__6144 (
            .O(N__31753),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__6143 (
            .O(N__31750),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__6142 (
            .O(N__31743),
            .I(N__31740));
    LocalMux I__6141 (
            .O(N__31740),
            .I(N__31736));
    CascadeMux I__6140 (
            .O(N__31739),
            .I(N__31733));
    Span4Mux_v I__6139 (
            .O(N__31736),
            .I(N__31730));
    InMux I__6138 (
            .O(N__31733),
            .I(N__31727));
    Span4Mux_v I__6137 (
            .O(N__31730),
            .I(N__31723));
    LocalMux I__6136 (
            .O(N__31727),
            .I(N__31719));
    CascadeMux I__6135 (
            .O(N__31726),
            .I(N__31716));
    Span4Mux_v I__6134 (
            .O(N__31723),
            .I(N__31713));
    InMux I__6133 (
            .O(N__31722),
            .I(N__31710));
    Span4Mux_h I__6132 (
            .O(N__31719),
            .I(N__31707));
    InMux I__6131 (
            .O(N__31716),
            .I(N__31704));
    Span4Mux_v I__6130 (
            .O(N__31713),
            .I(N__31699));
    LocalMux I__6129 (
            .O(N__31710),
            .I(N__31699));
    Span4Mux_v I__6128 (
            .O(N__31707),
            .I(N__31692));
    LocalMux I__6127 (
            .O(N__31704),
            .I(N__31692));
    Span4Mux_h I__6126 (
            .O(N__31699),
            .I(N__31692));
    Odrv4 I__6125 (
            .O(N__31692),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__6124 (
            .O(N__31689),
            .I(N__31686));
    LocalMux I__6123 (
            .O(N__31686),
            .I(N__31683));
    Odrv4 I__6122 (
            .O(N__31683),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__6121 (
            .O(N__31680),
            .I(N__31676));
    InMux I__6120 (
            .O(N__31679),
            .I(N__31673));
    LocalMux I__6119 (
            .O(N__31676),
            .I(N__31669));
    LocalMux I__6118 (
            .O(N__31673),
            .I(N__31666));
    InMux I__6117 (
            .O(N__31672),
            .I(N__31663));
    Span4Mux_v I__6116 (
            .O(N__31669),
            .I(N__31658));
    Span4Mux_v I__6115 (
            .O(N__31666),
            .I(N__31658));
    LocalMux I__6114 (
            .O(N__31663),
            .I(N__31654));
    Span4Mux_h I__6113 (
            .O(N__31658),
            .I(N__31651));
    InMux I__6112 (
            .O(N__31657),
            .I(N__31648));
    Odrv4 I__6111 (
            .O(N__31654),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__6110 (
            .O(N__31651),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__6109 (
            .O(N__31648),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__6108 (
            .O(N__31641),
            .I(N__31638));
    LocalMux I__6107 (
            .O(N__31638),
            .I(N__31635));
    Span4Mux_v I__6106 (
            .O(N__31635),
            .I(N__31630));
    InMux I__6105 (
            .O(N__31634),
            .I(N__31625));
    InMux I__6104 (
            .O(N__31633),
            .I(N__31625));
    Sp12to4 I__6103 (
            .O(N__31630),
            .I(N__31619));
    LocalMux I__6102 (
            .O(N__31625),
            .I(N__31619));
    InMux I__6101 (
            .O(N__31624),
            .I(N__31616));
    Odrv12 I__6100 (
            .O(N__31619),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__6099 (
            .O(N__31616),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__6098 (
            .O(N__31611),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__6097 (
            .O(N__31608),
            .I(N__31604));
    InMux I__6096 (
            .O(N__31607),
            .I(N__31601));
    LocalMux I__6095 (
            .O(N__31604),
            .I(N__31597));
    LocalMux I__6094 (
            .O(N__31601),
            .I(N__31594));
    InMux I__6093 (
            .O(N__31600),
            .I(N__31591));
    Span4Mux_h I__6092 (
            .O(N__31597),
            .I(N__31587));
    Span4Mux_v I__6091 (
            .O(N__31594),
            .I(N__31584));
    LocalMux I__6090 (
            .O(N__31591),
            .I(N__31581));
    InMux I__6089 (
            .O(N__31590),
            .I(N__31578));
    Odrv4 I__6088 (
            .O(N__31587),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__6087 (
            .O(N__31584),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv12 I__6086 (
            .O(N__31581),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__6085 (
            .O(N__31578),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__6084 (
            .O(N__31569),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__6083 (
            .O(N__31566),
            .I(N__31563));
    LocalMux I__6082 (
            .O(N__31563),
            .I(N__31559));
    InMux I__6081 (
            .O(N__31562),
            .I(N__31556));
    Span4Mux_v I__6080 (
            .O(N__31559),
            .I(N__31551));
    LocalMux I__6079 (
            .O(N__31556),
            .I(N__31551));
    Span4Mux_h I__6078 (
            .O(N__31551),
            .I(N__31546));
    InMux I__6077 (
            .O(N__31550),
            .I(N__31541));
    InMux I__6076 (
            .O(N__31549),
            .I(N__31541));
    Odrv4 I__6075 (
            .O(N__31546),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__6074 (
            .O(N__31541),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__6073 (
            .O(N__31536),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__6072 (
            .O(N__31533),
            .I(N__31530));
    LocalMux I__6071 (
            .O(N__31530),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ));
    InMux I__6070 (
            .O(N__31527),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__6069 (
            .O(N__31524),
            .I(N__31521));
    InMux I__6068 (
            .O(N__31521),
            .I(N__31518));
    LocalMux I__6067 (
            .O(N__31518),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__6066 (
            .O(N__31515),
            .I(N__31512));
    InMux I__6065 (
            .O(N__31512),
            .I(N__31509));
    LocalMux I__6064 (
            .O(N__31509),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__6063 (
            .O(N__31506),
            .I(N__31503));
    InMux I__6062 (
            .O(N__31503),
            .I(N__31500));
    LocalMux I__6061 (
            .O(N__31500),
            .I(N__31497));
    Odrv4 I__6060 (
            .O(N__31497),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__6059 (
            .O(N__31494),
            .I(N__31491));
    InMux I__6058 (
            .O(N__31491),
            .I(N__31488));
    LocalMux I__6057 (
            .O(N__31488),
            .I(N__31485));
    Odrv4 I__6056 (
            .O(N__31485),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__6055 (
            .O(N__31482),
            .I(N__31471));
    InMux I__6054 (
            .O(N__31481),
            .I(N__31471));
    InMux I__6053 (
            .O(N__31480),
            .I(N__31471));
    InMux I__6052 (
            .O(N__31479),
            .I(N__31466));
    InMux I__6051 (
            .O(N__31478),
            .I(N__31466));
    LocalMux I__6050 (
            .O(N__31471),
            .I(N__31456));
    LocalMux I__6049 (
            .O(N__31466),
            .I(N__31456));
    InMux I__6048 (
            .O(N__31465),
            .I(N__31453));
    InMux I__6047 (
            .O(N__31464),
            .I(N__31450));
    InMux I__6046 (
            .O(N__31463),
            .I(N__31447));
    InMux I__6045 (
            .O(N__31462),
            .I(N__31442));
    InMux I__6044 (
            .O(N__31461),
            .I(N__31442));
    Span12Mux_h I__6043 (
            .O(N__31456),
            .I(N__31439));
    LocalMux I__6042 (
            .O(N__31453),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__6041 (
            .O(N__31450),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__6040 (
            .O(N__31447),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    LocalMux I__6039 (
            .O(N__31442),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    Odrv12 I__6038 (
            .O(N__31439),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ));
    CascadeMux I__6037 (
            .O(N__31428),
            .I(N__31425));
    InMux I__6036 (
            .O(N__31425),
            .I(N__31422));
    LocalMux I__6035 (
            .O(N__31422),
            .I(N__31419));
    Odrv4 I__6034 (
            .O(N__31419),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__6033 (
            .O(N__31416),
            .I(N__31413));
    LocalMux I__6032 (
            .O(N__31413),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__6031 (
            .O(N__31410),
            .I(N__31407));
    InMux I__6030 (
            .O(N__31407),
            .I(N__31404));
    LocalMux I__6029 (
            .O(N__31404),
            .I(N__31401));
    Odrv4 I__6028 (
            .O(N__31401),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    InMux I__6027 (
            .O(N__31398),
            .I(N__31395));
    LocalMux I__6026 (
            .O(N__31395),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__6025 (
            .O(N__31392),
            .I(N__31389));
    InMux I__6024 (
            .O(N__31389),
            .I(N__31386));
    LocalMux I__6023 (
            .O(N__31386),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__6022 (
            .O(N__31383),
            .I(N__31380));
    LocalMux I__6021 (
            .O(N__31380),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__6020 (
            .O(N__31377),
            .I(N__31374));
    InMux I__6019 (
            .O(N__31374),
            .I(N__31371));
    LocalMux I__6018 (
            .O(N__31371),
            .I(N__31368));
    Odrv4 I__6017 (
            .O(N__31368),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__6016 (
            .O(N__31365),
            .I(N__31362));
    LocalMux I__6015 (
            .O(N__31362),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__6014 (
            .O(N__31359),
            .I(N__31356));
    InMux I__6013 (
            .O(N__31356),
            .I(N__31353));
    LocalMux I__6012 (
            .O(N__31353),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__6011 (
            .O(N__31350),
            .I(N__31347));
    LocalMux I__6010 (
            .O(N__31347),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__6009 (
            .O(N__31344),
            .I(N__31341));
    LocalMux I__6008 (
            .O(N__31341),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ));
    CascadeMux I__6007 (
            .O(N__31338),
            .I(N__31335));
    InMux I__6006 (
            .O(N__31335),
            .I(N__31332));
    LocalMux I__6005 (
            .O(N__31332),
            .I(N__31329));
    Odrv4 I__6004 (
            .O(N__31329),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__6003 (
            .O(N__31326),
            .I(N__31323));
    LocalMux I__6002 (
            .O(N__31323),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ));
    InMux I__6001 (
            .O(N__31320),
            .I(N__31317));
    LocalMux I__6000 (
            .O(N__31317),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ));
    CascadeMux I__5999 (
            .O(N__31314),
            .I(N__31311));
    InMux I__5998 (
            .O(N__31311),
            .I(N__31308));
    LocalMux I__5997 (
            .O(N__31308),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    InMux I__5996 (
            .O(N__31305),
            .I(N__31302));
    LocalMux I__5995 (
            .O(N__31302),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__5994 (
            .O(N__31299),
            .I(N__31296));
    InMux I__5993 (
            .O(N__31296),
            .I(N__31293));
    LocalMux I__5992 (
            .O(N__31293),
            .I(N__31290));
    Odrv4 I__5991 (
            .O(N__31290),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__5990 (
            .O(N__31287),
            .I(N__31284));
    LocalMux I__5989 (
            .O(N__31284),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__5988 (
            .O(N__31281),
            .I(N__31278));
    InMux I__5987 (
            .O(N__31278),
            .I(N__31275));
    LocalMux I__5986 (
            .O(N__31275),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    InMux I__5985 (
            .O(N__31272),
            .I(N__31269));
    LocalMux I__5984 (
            .O(N__31269),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__5983 (
            .O(N__31266),
            .I(N__31263));
    InMux I__5982 (
            .O(N__31263),
            .I(N__31260));
    LocalMux I__5981 (
            .O(N__31260),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__5980 (
            .O(N__31257),
            .I(N__31254));
    LocalMux I__5979 (
            .O(N__31254),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__5978 (
            .O(N__31251),
            .I(N__31248));
    InMux I__5977 (
            .O(N__31248),
            .I(N__31245));
    LocalMux I__5976 (
            .O(N__31245),
            .I(N__31242));
    Odrv4 I__5975 (
            .O(N__31242),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__5974 (
            .O(N__31239),
            .I(N__31236));
    LocalMux I__5973 (
            .O(N__31236),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__5972 (
            .O(N__31233),
            .I(N__31230));
    InMux I__5971 (
            .O(N__31230),
            .I(N__31227));
    LocalMux I__5970 (
            .O(N__31227),
            .I(N__31224));
    Span4Mux_h I__5969 (
            .O(N__31224),
            .I(N__31221));
    Odrv4 I__5968 (
            .O(N__31221),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__5967 (
            .O(N__31218),
            .I(N__31215));
    LocalMux I__5966 (
            .O(N__31215),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__5965 (
            .O(N__31212),
            .I(N__31209));
    LocalMux I__5964 (
            .O(N__31209),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__5963 (
            .O(N__31206),
            .I(N__31203));
    InMux I__5962 (
            .O(N__31203),
            .I(N__31200));
    LocalMux I__5961 (
            .O(N__31200),
            .I(N__31197));
    Odrv4 I__5960 (
            .O(N__31197),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__5959 (
            .O(N__31194),
            .I(N__31191));
    LocalMux I__5958 (
            .O(N__31191),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__5957 (
            .O(N__31188),
            .I(N__31183));
    InMux I__5956 (
            .O(N__31187),
            .I(N__31179));
    InMux I__5955 (
            .O(N__31186),
            .I(N__31176));
    InMux I__5954 (
            .O(N__31183),
            .I(N__31171));
    InMux I__5953 (
            .O(N__31182),
            .I(N__31171));
    LocalMux I__5952 (
            .O(N__31179),
            .I(N__31168));
    LocalMux I__5951 (
            .O(N__31176),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__5950 (
            .O(N__31171),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__5949 (
            .O(N__31168),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__5948 (
            .O(N__31161),
            .I(N__31155));
    InMux I__5947 (
            .O(N__31160),
            .I(N__31152));
    InMux I__5946 (
            .O(N__31159),
            .I(N__31147));
    InMux I__5945 (
            .O(N__31158),
            .I(N__31147));
    LocalMux I__5944 (
            .O(N__31155),
            .I(N__31144));
    LocalMux I__5943 (
            .O(N__31152),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__5942 (
            .O(N__31147),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__5941 (
            .O(N__31144),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__5940 (
            .O(N__31137),
            .I(N__31132));
    InMux I__5939 (
            .O(N__31136),
            .I(N__31128));
    InMux I__5938 (
            .O(N__31135),
            .I(N__31125));
    LocalMux I__5937 (
            .O(N__31132),
            .I(N__31122));
    InMux I__5936 (
            .O(N__31131),
            .I(N__31119));
    LocalMux I__5935 (
            .O(N__31128),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__5934 (
            .O(N__31125),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv12 I__5933 (
            .O(N__31122),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__5932 (
            .O(N__31119),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__5931 (
            .O(N__31110),
            .I(N__31107));
    LocalMux I__5930 (
            .O(N__31107),
            .I(N__31104));
    Span4Mux_s2_v I__5929 (
            .O(N__31104),
            .I(N__31101));
    Span4Mux_v I__5928 (
            .O(N__31101),
            .I(N__31098));
    Odrv4 I__5927 (
            .O(N__31098),
            .I(\current_shift_inst.timer_s1.N_185_i ));
    InMux I__5926 (
            .O(N__31095),
            .I(N__31090));
    InMux I__5925 (
            .O(N__31094),
            .I(N__31087));
    InMux I__5924 (
            .O(N__31093),
            .I(N__31084));
    LocalMux I__5923 (
            .O(N__31090),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__5922 (
            .O(N__31087),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    LocalMux I__5921 (
            .O(N__31084),
            .I(\delay_measurement_inst.prev_tr_sigZ0 ));
    InMux I__5920 (
            .O(N__31077),
            .I(N__31072));
    InMux I__5919 (
            .O(N__31076),
            .I(N__31069));
    InMux I__5918 (
            .O(N__31075),
            .I(N__31066));
    LocalMux I__5917 (
            .O(N__31072),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__5916 (
            .O(N__31069),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    LocalMux I__5915 (
            .O(N__31066),
            .I(\delay_measurement_inst.tr_stateZ0Z_0 ));
    InMux I__5914 (
            .O(N__31059),
            .I(N__31056));
    LocalMux I__5913 (
            .O(N__31056),
            .I(N__31053));
    Span4Mux_h I__5912 (
            .O(N__31053),
            .I(N__31050));
    Sp12to4 I__5911 (
            .O(N__31050),
            .I(N__31047));
    Odrv12 I__5910 (
            .O(N__31047),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    InMux I__5909 (
            .O(N__31044),
            .I(N__31041));
    LocalMux I__5908 (
            .O(N__31041),
            .I(\phase_controller_inst2.start_timer_hc_RNO_0_0 ));
    InMux I__5907 (
            .O(N__31038),
            .I(N__31035));
    LocalMux I__5906 (
            .O(N__31035),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__5905 (
            .O(N__31032),
            .I(N__31029));
    InMux I__5904 (
            .O(N__31029),
            .I(N__31026));
    LocalMux I__5903 (
            .O(N__31026),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__5902 (
            .O(N__31023),
            .I(N__31020));
    InMux I__5901 (
            .O(N__31020),
            .I(N__31017));
    LocalMux I__5900 (
            .O(N__31017),
            .I(N__31014));
    Odrv4 I__5899 (
            .O(N__31014),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__5898 (
            .O(N__31011),
            .I(N__31008));
    LocalMux I__5897 (
            .O(N__31008),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__5896 (
            .O(N__31005),
            .I(N__31002));
    InMux I__5895 (
            .O(N__31002),
            .I(N__30999));
    LocalMux I__5894 (
            .O(N__30999),
            .I(N__30996));
    Odrv4 I__5893 (
            .O(N__30996),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__5892 (
            .O(N__30993),
            .I(N__30990));
    LocalMux I__5891 (
            .O(N__30990),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__5890 (
            .O(N__30987),
            .I(N__30984));
    LocalMux I__5889 (
            .O(N__30984),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__5888 (
            .O(N__30981),
            .I(N__30978));
    LocalMux I__5887 (
            .O(N__30978),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__5886 (
            .O(N__30975),
            .I(N__30972));
    LocalMux I__5885 (
            .O(N__30972),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__5884 (
            .O(N__30969),
            .I(N__30965));
    InMux I__5883 (
            .O(N__30968),
            .I(N__30962));
    LocalMux I__5882 (
            .O(N__30965),
            .I(N__30959));
    LocalMux I__5881 (
            .O(N__30962),
            .I(N__30956));
    Span4Mux_h I__5880 (
            .O(N__30959),
            .I(N__30953));
    Odrv12 I__5879 (
            .O(N__30956),
            .I(state_ns_i_a3_1));
    Odrv4 I__5878 (
            .O(N__30953),
            .I(state_ns_i_a3_1));
    InMux I__5877 (
            .O(N__30948),
            .I(N__30939));
    InMux I__5876 (
            .O(N__30947),
            .I(N__30932));
    InMux I__5875 (
            .O(N__30946),
            .I(N__30932));
    InMux I__5874 (
            .O(N__30945),
            .I(N__30932));
    InMux I__5873 (
            .O(N__30944),
            .I(N__30927));
    InMux I__5872 (
            .O(N__30943),
            .I(N__30927));
    CascadeMux I__5871 (
            .O(N__30942),
            .I(N__30912));
    LocalMux I__5870 (
            .O(N__30939),
            .I(N__30904));
    LocalMux I__5869 (
            .O(N__30932),
            .I(N__30899));
    LocalMux I__5868 (
            .O(N__30927),
            .I(N__30899));
    InMux I__5867 (
            .O(N__30926),
            .I(N__30884));
    InMux I__5866 (
            .O(N__30925),
            .I(N__30884));
    InMux I__5865 (
            .O(N__30924),
            .I(N__30884));
    InMux I__5864 (
            .O(N__30923),
            .I(N__30884));
    InMux I__5863 (
            .O(N__30922),
            .I(N__30884));
    InMux I__5862 (
            .O(N__30921),
            .I(N__30884));
    InMux I__5861 (
            .O(N__30920),
            .I(N__30884));
    InMux I__5860 (
            .O(N__30919),
            .I(N__30871));
    InMux I__5859 (
            .O(N__30918),
            .I(N__30871));
    InMux I__5858 (
            .O(N__30917),
            .I(N__30871));
    InMux I__5857 (
            .O(N__30916),
            .I(N__30871));
    InMux I__5856 (
            .O(N__30915),
            .I(N__30871));
    InMux I__5855 (
            .O(N__30912),
            .I(N__30871));
    InMux I__5854 (
            .O(N__30911),
            .I(N__30860));
    InMux I__5853 (
            .O(N__30910),
            .I(N__30860));
    InMux I__5852 (
            .O(N__30909),
            .I(N__30860));
    InMux I__5851 (
            .O(N__30908),
            .I(N__30860));
    InMux I__5850 (
            .O(N__30907),
            .I(N__30860));
    Span4Mux_v I__5849 (
            .O(N__30904),
            .I(N__30856));
    Span4Mux_v I__5848 (
            .O(N__30899),
            .I(N__30853));
    LocalMux I__5847 (
            .O(N__30884),
            .I(N__30846));
    LocalMux I__5846 (
            .O(N__30871),
            .I(N__30846));
    LocalMux I__5845 (
            .O(N__30860),
            .I(N__30846));
    InMux I__5844 (
            .O(N__30859),
            .I(N__30843));
    Odrv4 I__5843 (
            .O(N__30856),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__5842 (
            .O(N__30853),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__5841 (
            .O(N__30846),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__5840 (
            .O(N__30843),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    InMux I__5839 (
            .O(N__30834),
            .I(N__30831));
    LocalMux I__5838 (
            .O(N__30831),
            .I(N__30826));
    InMux I__5837 (
            .O(N__30830),
            .I(N__30823));
    InMux I__5836 (
            .O(N__30829),
            .I(N__30820));
    Span4Mux_v I__5835 (
            .O(N__30826),
            .I(N__30817));
    LocalMux I__5834 (
            .O(N__30823),
            .I(N__30812));
    LocalMux I__5833 (
            .O(N__30820),
            .I(N__30812));
    Odrv4 I__5832 (
            .O(N__30817),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__5831 (
            .O(N__30812),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__5830 (
            .O(N__30807),
            .I(N__30804));
    LocalMux I__5829 (
            .O(N__30804),
            .I(N__30801));
    Span4Mux_h I__5828 (
            .O(N__30801),
            .I(N__30798));
    Odrv4 I__5827 (
            .O(N__30798),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__5826 (
            .O(N__30795),
            .I(N__30792));
    LocalMux I__5825 (
            .O(N__30792),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__5824 (
            .O(N__30789),
            .I(N__30786));
    LocalMux I__5823 (
            .O(N__30786),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__5822 (
            .O(N__30783),
            .I(N__30780));
    LocalMux I__5821 (
            .O(N__30780),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__5820 (
            .O(N__30777),
            .I(N__30774));
    LocalMux I__5819 (
            .O(N__30774),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__5818 (
            .O(N__30771),
            .I(N__30768));
    LocalMux I__5817 (
            .O(N__30768),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__5816 (
            .O(N__30765),
            .I(N__30762));
    LocalMux I__5815 (
            .O(N__30762),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__5814 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__5813 (
            .O(N__30756),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__5812 (
            .O(N__30753),
            .I(N__30750));
    LocalMux I__5811 (
            .O(N__30750),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__5810 (
            .O(N__30747),
            .I(N__30744));
    LocalMux I__5809 (
            .O(N__30744),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__5808 (
            .O(N__30741),
            .I(N__30738));
    LocalMux I__5807 (
            .O(N__30738),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__5806 (
            .O(N__30735),
            .I(N__30732));
    LocalMux I__5805 (
            .O(N__30732),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__5804 (
            .O(N__30729),
            .I(N__30726));
    LocalMux I__5803 (
            .O(N__30726),
            .I(N__30723));
    Span4Mux_h I__5802 (
            .O(N__30723),
            .I(N__30718));
    InMux I__5801 (
            .O(N__30722),
            .I(N__30715));
    InMux I__5800 (
            .O(N__30721),
            .I(N__30712));
    Odrv4 I__5799 (
            .O(N__30718),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__5798 (
            .O(N__30715),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__5797 (
            .O(N__30712),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__5796 (
            .O(N__30705),
            .I(N__30702));
    LocalMux I__5795 (
            .O(N__30702),
            .I(N__30699));
    Span4Mux_v I__5794 (
            .O(N__30699),
            .I(N__30696));
    Odrv4 I__5793 (
            .O(N__30696),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    CascadeMux I__5792 (
            .O(N__30693),
            .I(N__30683));
    CascadeMux I__5791 (
            .O(N__30692),
            .I(N__30680));
    CascadeMux I__5790 (
            .O(N__30691),
            .I(N__30661));
    CascadeMux I__5789 (
            .O(N__30690),
            .I(N__30658));
    CascadeMux I__5788 (
            .O(N__30689),
            .I(N__30655));
    CascadeMux I__5787 (
            .O(N__30688),
            .I(N__30652));
    CascadeMux I__5786 (
            .O(N__30687),
            .I(N__30649));
    CascadeMux I__5785 (
            .O(N__30686),
            .I(N__30644));
    InMux I__5784 (
            .O(N__30683),
            .I(N__30641));
    InMux I__5783 (
            .O(N__30680),
            .I(N__30638));
    InMux I__5782 (
            .O(N__30679),
            .I(N__30635));
    CascadeMux I__5781 (
            .O(N__30678),
            .I(N__30632));
    CascadeMux I__5780 (
            .O(N__30677),
            .I(N__30629));
    CascadeMux I__5779 (
            .O(N__30676),
            .I(N__30626));
    CascadeMux I__5778 (
            .O(N__30675),
            .I(N__30616));
    CascadeMux I__5777 (
            .O(N__30674),
            .I(N__30611));
    InMux I__5776 (
            .O(N__30673),
            .I(N__30607));
    CascadeMux I__5775 (
            .O(N__30672),
            .I(N__30599));
    CascadeMux I__5774 (
            .O(N__30671),
            .I(N__30592));
    CascadeMux I__5773 (
            .O(N__30670),
            .I(N__30589));
    CascadeMux I__5772 (
            .O(N__30669),
            .I(N__30585));
    CascadeMux I__5771 (
            .O(N__30668),
            .I(N__30582));
    CascadeMux I__5770 (
            .O(N__30667),
            .I(N__30579));
    CascadeMux I__5769 (
            .O(N__30666),
            .I(N__30576));
    CascadeMux I__5768 (
            .O(N__30665),
            .I(N__30573));
    CascadeMux I__5767 (
            .O(N__30664),
            .I(N__30570));
    InMux I__5766 (
            .O(N__30661),
            .I(N__30563));
    InMux I__5765 (
            .O(N__30658),
            .I(N__30560));
    InMux I__5764 (
            .O(N__30655),
            .I(N__30555));
    InMux I__5763 (
            .O(N__30652),
            .I(N__30555));
    InMux I__5762 (
            .O(N__30649),
            .I(N__30548));
    InMux I__5761 (
            .O(N__30648),
            .I(N__30548));
    InMux I__5760 (
            .O(N__30647),
            .I(N__30548));
    InMux I__5759 (
            .O(N__30644),
            .I(N__30545));
    LocalMux I__5758 (
            .O(N__30641),
            .I(N__30538));
    LocalMux I__5757 (
            .O(N__30638),
            .I(N__30538));
    LocalMux I__5756 (
            .O(N__30635),
            .I(N__30538));
    InMux I__5755 (
            .O(N__30632),
            .I(N__30531));
    InMux I__5754 (
            .O(N__30629),
            .I(N__30531));
    InMux I__5753 (
            .O(N__30626),
            .I(N__30531));
    CascadeMux I__5752 (
            .O(N__30625),
            .I(N__30528));
    CascadeMux I__5751 (
            .O(N__30624),
            .I(N__30525));
    CascadeMux I__5750 (
            .O(N__30623),
            .I(N__30522));
    CascadeMux I__5749 (
            .O(N__30622),
            .I(N__30519));
    CascadeMux I__5748 (
            .O(N__30621),
            .I(N__30516));
    CascadeMux I__5747 (
            .O(N__30620),
            .I(N__30513));
    CascadeMux I__5746 (
            .O(N__30619),
            .I(N__30510));
    InMux I__5745 (
            .O(N__30616),
            .I(N__30507));
    InMux I__5744 (
            .O(N__30615),
            .I(N__30504));
    InMux I__5743 (
            .O(N__30614),
            .I(N__30501));
    InMux I__5742 (
            .O(N__30611),
            .I(N__30498));
    CascadeMux I__5741 (
            .O(N__30610),
            .I(N__30495));
    LocalMux I__5740 (
            .O(N__30607),
            .I(N__30489));
    CascadeMux I__5739 (
            .O(N__30606),
            .I(N__30486));
    CascadeMux I__5738 (
            .O(N__30605),
            .I(N__30483));
    CascadeMux I__5737 (
            .O(N__30604),
            .I(N__30479));
    CascadeMux I__5736 (
            .O(N__30603),
            .I(N__30476));
    CascadeMux I__5735 (
            .O(N__30602),
            .I(N__30472));
    InMux I__5734 (
            .O(N__30599),
            .I(N__30461));
    CascadeMux I__5733 (
            .O(N__30598),
            .I(N__30455));
    CascadeMux I__5732 (
            .O(N__30597),
            .I(N__30452));
    CascadeMux I__5731 (
            .O(N__30596),
            .I(N__30449));
    CascadeMux I__5730 (
            .O(N__30595),
            .I(N__30445));
    InMux I__5729 (
            .O(N__30592),
            .I(N__30421));
    InMux I__5728 (
            .O(N__30589),
            .I(N__30412));
    InMux I__5727 (
            .O(N__30588),
            .I(N__30412));
    InMux I__5726 (
            .O(N__30585),
            .I(N__30412));
    InMux I__5725 (
            .O(N__30582),
            .I(N__30412));
    InMux I__5724 (
            .O(N__30579),
            .I(N__30403));
    InMux I__5723 (
            .O(N__30576),
            .I(N__30403));
    InMux I__5722 (
            .O(N__30573),
            .I(N__30403));
    InMux I__5721 (
            .O(N__30570),
            .I(N__30403));
    CascadeMux I__5720 (
            .O(N__30569),
            .I(N__30400));
    CascadeMux I__5719 (
            .O(N__30568),
            .I(N__30397));
    CascadeMux I__5718 (
            .O(N__30567),
            .I(N__30394));
    CascadeMux I__5717 (
            .O(N__30566),
            .I(N__30390));
    LocalMux I__5716 (
            .O(N__30563),
            .I(N__30375));
    LocalMux I__5715 (
            .O(N__30560),
            .I(N__30375));
    LocalMux I__5714 (
            .O(N__30555),
            .I(N__30375));
    LocalMux I__5713 (
            .O(N__30548),
            .I(N__30375));
    LocalMux I__5712 (
            .O(N__30545),
            .I(N__30375));
    Span4Mux_v I__5711 (
            .O(N__30538),
            .I(N__30375));
    LocalMux I__5710 (
            .O(N__30531),
            .I(N__30375));
    InMux I__5709 (
            .O(N__30528),
            .I(N__30366));
    InMux I__5708 (
            .O(N__30525),
            .I(N__30366));
    InMux I__5707 (
            .O(N__30522),
            .I(N__30366));
    InMux I__5706 (
            .O(N__30519),
            .I(N__30366));
    InMux I__5705 (
            .O(N__30516),
            .I(N__30359));
    InMux I__5704 (
            .O(N__30513),
            .I(N__30359));
    InMux I__5703 (
            .O(N__30510),
            .I(N__30359));
    LocalMux I__5702 (
            .O(N__30507),
            .I(N__30354));
    LocalMux I__5701 (
            .O(N__30504),
            .I(N__30354));
    LocalMux I__5700 (
            .O(N__30501),
            .I(N__30351));
    LocalMux I__5699 (
            .O(N__30498),
            .I(N__30343));
    InMux I__5698 (
            .O(N__30495),
            .I(N__30338));
    InMux I__5697 (
            .O(N__30494),
            .I(N__30338));
    CascadeMux I__5696 (
            .O(N__30493),
            .I(N__30335));
    CascadeMux I__5695 (
            .O(N__30492),
            .I(N__30329));
    Span4Mux_h I__5694 (
            .O(N__30489),
            .I(N__30326));
    InMux I__5693 (
            .O(N__30486),
            .I(N__30323));
    InMux I__5692 (
            .O(N__30483),
            .I(N__30316));
    InMux I__5691 (
            .O(N__30482),
            .I(N__30316));
    InMux I__5690 (
            .O(N__30479),
            .I(N__30316));
    InMux I__5689 (
            .O(N__30476),
            .I(N__30309));
    InMux I__5688 (
            .O(N__30475),
            .I(N__30309));
    InMux I__5687 (
            .O(N__30472),
            .I(N__30309));
    InMux I__5686 (
            .O(N__30471),
            .I(N__30304));
    InMux I__5685 (
            .O(N__30470),
            .I(N__30304));
    CascadeMux I__5684 (
            .O(N__30469),
            .I(N__30301));
    CascadeMux I__5683 (
            .O(N__30468),
            .I(N__30298));
    CascadeMux I__5682 (
            .O(N__30467),
            .I(N__30295));
    CascadeMux I__5681 (
            .O(N__30466),
            .I(N__30292));
    CascadeMux I__5680 (
            .O(N__30465),
            .I(N__30289));
    CascadeMux I__5679 (
            .O(N__30464),
            .I(N__30286));
    LocalMux I__5678 (
            .O(N__30461),
            .I(N__30269));
    CascadeMux I__5677 (
            .O(N__30460),
            .I(N__30265));
    CascadeMux I__5676 (
            .O(N__30459),
            .I(N__30262));
    CascadeMux I__5675 (
            .O(N__30458),
            .I(N__30259));
    InMux I__5674 (
            .O(N__30455),
            .I(N__30248));
    InMux I__5673 (
            .O(N__30452),
            .I(N__30248));
    InMux I__5672 (
            .O(N__30449),
            .I(N__30248));
    InMux I__5671 (
            .O(N__30448),
            .I(N__30248));
    InMux I__5670 (
            .O(N__30445),
            .I(N__30248));
    CascadeMux I__5669 (
            .O(N__30444),
            .I(N__30245));
    CascadeMux I__5668 (
            .O(N__30443),
            .I(N__30242));
    CascadeMux I__5667 (
            .O(N__30442),
            .I(N__30239));
    CascadeMux I__5666 (
            .O(N__30441),
            .I(N__30235));
    CascadeMux I__5665 (
            .O(N__30440),
            .I(N__30232));
    CascadeMux I__5664 (
            .O(N__30439),
            .I(N__30229));
    CascadeMux I__5663 (
            .O(N__30438),
            .I(N__30226));
    CascadeMux I__5662 (
            .O(N__30437),
            .I(N__30223));
    CascadeMux I__5661 (
            .O(N__30436),
            .I(N__30220));
    CascadeMux I__5660 (
            .O(N__30435),
            .I(N__30217));
    CascadeMux I__5659 (
            .O(N__30434),
            .I(N__30214));
    CascadeMux I__5658 (
            .O(N__30433),
            .I(N__30211));
    CascadeMux I__5657 (
            .O(N__30432),
            .I(N__30208));
    CascadeMux I__5656 (
            .O(N__30431),
            .I(N__30205));
    CascadeMux I__5655 (
            .O(N__30430),
            .I(N__30202));
    CascadeMux I__5654 (
            .O(N__30429),
            .I(N__30199));
    CascadeMux I__5653 (
            .O(N__30428),
            .I(N__30196));
    CascadeMux I__5652 (
            .O(N__30427),
            .I(N__30193));
    CascadeMux I__5651 (
            .O(N__30426),
            .I(N__30190));
    CascadeMux I__5650 (
            .O(N__30425),
            .I(N__30187));
    CascadeMux I__5649 (
            .O(N__30424),
            .I(N__30183));
    LocalMux I__5648 (
            .O(N__30421),
            .I(N__30176));
    LocalMux I__5647 (
            .O(N__30412),
            .I(N__30176));
    LocalMux I__5646 (
            .O(N__30403),
            .I(N__30176));
    InMux I__5645 (
            .O(N__30400),
            .I(N__30171));
    InMux I__5644 (
            .O(N__30397),
            .I(N__30171));
    InMux I__5643 (
            .O(N__30394),
            .I(N__30164));
    InMux I__5642 (
            .O(N__30393),
            .I(N__30164));
    InMux I__5641 (
            .O(N__30390),
            .I(N__30164));
    Span4Mux_v I__5640 (
            .O(N__30375),
            .I(N__30157));
    LocalMux I__5639 (
            .O(N__30366),
            .I(N__30157));
    LocalMux I__5638 (
            .O(N__30359),
            .I(N__30157));
    Span4Mux_h I__5637 (
            .O(N__30354),
            .I(N__30152));
    Span4Mux_v I__5636 (
            .O(N__30351),
            .I(N__30152));
    CascadeMux I__5635 (
            .O(N__30350),
            .I(N__30149));
    CascadeMux I__5634 (
            .O(N__30349),
            .I(N__30146));
    CascadeMux I__5633 (
            .O(N__30348),
            .I(N__30142));
    CascadeMux I__5632 (
            .O(N__30347),
            .I(N__30138));
    CascadeMux I__5631 (
            .O(N__30346),
            .I(N__30135));
    Span4Mux_v I__5630 (
            .O(N__30343),
            .I(N__30130));
    LocalMux I__5629 (
            .O(N__30338),
            .I(N__30130));
    InMux I__5628 (
            .O(N__30335),
            .I(N__30127));
    CascadeMux I__5627 (
            .O(N__30334),
            .I(N__30124));
    CascadeMux I__5626 (
            .O(N__30333),
            .I(N__30121));
    InMux I__5625 (
            .O(N__30332),
            .I(N__30118));
    InMux I__5624 (
            .O(N__30329),
            .I(N__30115));
    Span4Mux_v I__5623 (
            .O(N__30326),
            .I(N__30104));
    LocalMux I__5622 (
            .O(N__30323),
            .I(N__30104));
    LocalMux I__5621 (
            .O(N__30316),
            .I(N__30104));
    LocalMux I__5620 (
            .O(N__30309),
            .I(N__30104));
    LocalMux I__5619 (
            .O(N__30304),
            .I(N__30104));
    InMux I__5618 (
            .O(N__30301),
            .I(N__30099));
    InMux I__5617 (
            .O(N__30298),
            .I(N__30099));
    InMux I__5616 (
            .O(N__30295),
            .I(N__30090));
    InMux I__5615 (
            .O(N__30292),
            .I(N__30090));
    InMux I__5614 (
            .O(N__30289),
            .I(N__30090));
    InMux I__5613 (
            .O(N__30286),
            .I(N__30090));
    CascadeMux I__5612 (
            .O(N__30285),
            .I(N__30087));
    CascadeMux I__5611 (
            .O(N__30284),
            .I(N__30084));
    CascadeMux I__5610 (
            .O(N__30283),
            .I(N__30081));
    CascadeMux I__5609 (
            .O(N__30282),
            .I(N__30078));
    CascadeMux I__5608 (
            .O(N__30281),
            .I(N__30075));
    CascadeMux I__5607 (
            .O(N__30280),
            .I(N__30072));
    CascadeMux I__5606 (
            .O(N__30279),
            .I(N__30069));
    CascadeMux I__5605 (
            .O(N__30278),
            .I(N__30066));
    CascadeMux I__5604 (
            .O(N__30277),
            .I(N__30063));
    CascadeMux I__5603 (
            .O(N__30276),
            .I(N__30060));
    CascadeMux I__5602 (
            .O(N__30275),
            .I(N__30057));
    CascadeMux I__5601 (
            .O(N__30274),
            .I(N__30054));
    CascadeMux I__5600 (
            .O(N__30273),
            .I(N__30051));
    CascadeMux I__5599 (
            .O(N__30272),
            .I(N__30048));
    Span4Mux_v I__5598 (
            .O(N__30269),
            .I(N__30045));
    InMux I__5597 (
            .O(N__30268),
            .I(N__30036));
    InMux I__5596 (
            .O(N__30265),
            .I(N__30036));
    InMux I__5595 (
            .O(N__30262),
            .I(N__30036));
    InMux I__5594 (
            .O(N__30259),
            .I(N__30036));
    LocalMux I__5593 (
            .O(N__30248),
            .I(N__30033));
    InMux I__5592 (
            .O(N__30245),
            .I(N__30024));
    InMux I__5591 (
            .O(N__30242),
            .I(N__30024));
    InMux I__5590 (
            .O(N__30239),
            .I(N__30024));
    InMux I__5589 (
            .O(N__30238),
            .I(N__30024));
    InMux I__5588 (
            .O(N__30235),
            .I(N__30015));
    InMux I__5587 (
            .O(N__30232),
            .I(N__30015));
    InMux I__5586 (
            .O(N__30229),
            .I(N__30015));
    InMux I__5585 (
            .O(N__30226),
            .I(N__30015));
    InMux I__5584 (
            .O(N__30223),
            .I(N__30006));
    InMux I__5583 (
            .O(N__30220),
            .I(N__30006));
    InMux I__5582 (
            .O(N__30217),
            .I(N__30006));
    InMux I__5581 (
            .O(N__30214),
            .I(N__30006));
    InMux I__5580 (
            .O(N__30211),
            .I(N__29997));
    InMux I__5579 (
            .O(N__30208),
            .I(N__29997));
    InMux I__5578 (
            .O(N__30205),
            .I(N__29997));
    InMux I__5577 (
            .O(N__30202),
            .I(N__29997));
    InMux I__5576 (
            .O(N__30199),
            .I(N__29988));
    InMux I__5575 (
            .O(N__30196),
            .I(N__29988));
    InMux I__5574 (
            .O(N__30193),
            .I(N__29988));
    InMux I__5573 (
            .O(N__30190),
            .I(N__29988));
    InMux I__5572 (
            .O(N__30187),
            .I(N__29981));
    InMux I__5571 (
            .O(N__30186),
            .I(N__29981));
    InMux I__5570 (
            .O(N__30183),
            .I(N__29981));
    Span4Mux_v I__5569 (
            .O(N__30176),
            .I(N__29974));
    LocalMux I__5568 (
            .O(N__30171),
            .I(N__29974));
    LocalMux I__5567 (
            .O(N__30164),
            .I(N__29974));
    Span4Mux_h I__5566 (
            .O(N__30157),
            .I(N__29969));
    Span4Mux_h I__5565 (
            .O(N__30152),
            .I(N__29969));
    InMux I__5564 (
            .O(N__30149),
            .I(N__29960));
    InMux I__5563 (
            .O(N__30146),
            .I(N__29960));
    InMux I__5562 (
            .O(N__30145),
            .I(N__29960));
    InMux I__5561 (
            .O(N__30142),
            .I(N__29960));
    InMux I__5560 (
            .O(N__30141),
            .I(N__29953));
    InMux I__5559 (
            .O(N__30138),
            .I(N__29953));
    InMux I__5558 (
            .O(N__30135),
            .I(N__29953));
    Span4Mux_h I__5557 (
            .O(N__30130),
            .I(N__29948));
    LocalMux I__5556 (
            .O(N__30127),
            .I(N__29948));
    InMux I__5555 (
            .O(N__30124),
            .I(N__29945));
    InMux I__5554 (
            .O(N__30121),
            .I(N__29942));
    LocalMux I__5553 (
            .O(N__30118),
            .I(N__29937));
    LocalMux I__5552 (
            .O(N__30115),
            .I(N__29937));
    Span4Mux_h I__5551 (
            .O(N__30104),
            .I(N__29930));
    LocalMux I__5550 (
            .O(N__30099),
            .I(N__29930));
    LocalMux I__5549 (
            .O(N__30090),
            .I(N__29930));
    InMux I__5548 (
            .O(N__30087),
            .I(N__29921));
    InMux I__5547 (
            .O(N__30084),
            .I(N__29921));
    InMux I__5546 (
            .O(N__30081),
            .I(N__29921));
    InMux I__5545 (
            .O(N__30078),
            .I(N__29921));
    InMux I__5544 (
            .O(N__30075),
            .I(N__29912));
    InMux I__5543 (
            .O(N__30072),
            .I(N__29912));
    InMux I__5542 (
            .O(N__30069),
            .I(N__29912));
    InMux I__5541 (
            .O(N__30066),
            .I(N__29912));
    InMux I__5540 (
            .O(N__30063),
            .I(N__29903));
    InMux I__5539 (
            .O(N__30060),
            .I(N__29903));
    InMux I__5538 (
            .O(N__30057),
            .I(N__29903));
    InMux I__5537 (
            .O(N__30054),
            .I(N__29903));
    InMux I__5536 (
            .O(N__30051),
            .I(N__29898));
    InMux I__5535 (
            .O(N__30048),
            .I(N__29898));
    Span4Mux_v I__5534 (
            .O(N__30045),
            .I(N__29879));
    LocalMux I__5533 (
            .O(N__30036),
            .I(N__29879));
    Span4Mux_h I__5532 (
            .O(N__30033),
            .I(N__29879));
    LocalMux I__5531 (
            .O(N__30024),
            .I(N__29879));
    LocalMux I__5530 (
            .O(N__30015),
            .I(N__29879));
    LocalMux I__5529 (
            .O(N__30006),
            .I(N__29879));
    LocalMux I__5528 (
            .O(N__29997),
            .I(N__29879));
    LocalMux I__5527 (
            .O(N__29988),
            .I(N__29879));
    LocalMux I__5526 (
            .O(N__29981),
            .I(N__29879));
    Span4Mux_h I__5525 (
            .O(N__29974),
            .I(N__29870));
    Span4Mux_v I__5524 (
            .O(N__29969),
            .I(N__29870));
    LocalMux I__5523 (
            .O(N__29960),
            .I(N__29870));
    LocalMux I__5522 (
            .O(N__29953),
            .I(N__29870));
    Odrv4 I__5521 (
            .O(N__29948),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5520 (
            .O(N__29945),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5519 (
            .O(N__29942),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__5518 (
            .O(N__29937),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__5517 (
            .O(N__29930),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5516 (
            .O(N__29921),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5515 (
            .O(N__29912),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5514 (
            .O(N__29903),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5513 (
            .O(N__29898),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__5512 (
            .O(N__29879),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__5511 (
            .O(N__29870),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__5510 (
            .O(N__29847),
            .I(N__29838));
    CascadeMux I__5509 (
            .O(N__29846),
            .I(N__29829));
    InMux I__5508 (
            .O(N__29845),
            .I(N__29825));
    CascadeMux I__5507 (
            .O(N__29844),
            .I(N__29804));
    InMux I__5506 (
            .O(N__29843),
            .I(N__29796));
    InMux I__5505 (
            .O(N__29842),
            .I(N__29793));
    InMux I__5504 (
            .O(N__29841),
            .I(N__29784));
    InMux I__5503 (
            .O(N__29838),
            .I(N__29784));
    InMux I__5502 (
            .O(N__29837),
            .I(N__29784));
    InMux I__5501 (
            .O(N__29836),
            .I(N__29784));
    InMux I__5500 (
            .O(N__29835),
            .I(N__29777));
    InMux I__5499 (
            .O(N__29834),
            .I(N__29777));
    InMux I__5498 (
            .O(N__29833),
            .I(N__29768));
    InMux I__5497 (
            .O(N__29832),
            .I(N__29768));
    InMux I__5496 (
            .O(N__29829),
            .I(N__29768));
    InMux I__5495 (
            .O(N__29828),
            .I(N__29768));
    LocalMux I__5494 (
            .O(N__29825),
            .I(N__29764));
    InMux I__5493 (
            .O(N__29824),
            .I(N__29761));
    InMux I__5492 (
            .O(N__29823),
            .I(N__29756));
    InMux I__5491 (
            .O(N__29822),
            .I(N__29756));
    InMux I__5490 (
            .O(N__29821),
            .I(N__29747));
    InMux I__5489 (
            .O(N__29820),
            .I(N__29747));
    InMux I__5488 (
            .O(N__29819),
            .I(N__29747));
    InMux I__5487 (
            .O(N__29818),
            .I(N__29747));
    InMux I__5486 (
            .O(N__29817),
            .I(N__29740));
    InMux I__5485 (
            .O(N__29816),
            .I(N__29740));
    InMux I__5484 (
            .O(N__29815),
            .I(N__29740));
    InMux I__5483 (
            .O(N__29814),
            .I(N__29737));
    InMux I__5482 (
            .O(N__29813),
            .I(N__29722));
    InMux I__5481 (
            .O(N__29812),
            .I(N__29722));
    InMux I__5480 (
            .O(N__29811),
            .I(N__29722));
    InMux I__5479 (
            .O(N__29810),
            .I(N__29722));
    InMux I__5478 (
            .O(N__29809),
            .I(N__29719));
    InMux I__5477 (
            .O(N__29808),
            .I(N__29710));
    InMux I__5476 (
            .O(N__29807),
            .I(N__29710));
    InMux I__5475 (
            .O(N__29804),
            .I(N__29710));
    InMux I__5474 (
            .O(N__29803),
            .I(N__29710));
    InMux I__5473 (
            .O(N__29802),
            .I(N__29693));
    InMux I__5472 (
            .O(N__29801),
            .I(N__29687));
    InMux I__5471 (
            .O(N__29800),
            .I(N__29682));
    InMux I__5470 (
            .O(N__29799),
            .I(N__29682));
    LocalMux I__5469 (
            .O(N__29796),
            .I(N__29675));
    LocalMux I__5468 (
            .O(N__29793),
            .I(N__29675));
    LocalMux I__5467 (
            .O(N__29784),
            .I(N__29675));
    InMux I__5466 (
            .O(N__29783),
            .I(N__29670));
    InMux I__5465 (
            .O(N__29782),
            .I(N__29670));
    LocalMux I__5464 (
            .O(N__29777),
            .I(N__29665));
    LocalMux I__5463 (
            .O(N__29768),
            .I(N__29665));
    InMux I__5462 (
            .O(N__29767),
            .I(N__29662));
    Span4Mux_h I__5461 (
            .O(N__29764),
            .I(N__29651));
    LocalMux I__5460 (
            .O(N__29761),
            .I(N__29651));
    LocalMux I__5459 (
            .O(N__29756),
            .I(N__29651));
    LocalMux I__5458 (
            .O(N__29747),
            .I(N__29651));
    LocalMux I__5457 (
            .O(N__29740),
            .I(N__29651));
    LocalMux I__5456 (
            .O(N__29737),
            .I(N__29648));
    InMux I__5455 (
            .O(N__29736),
            .I(N__29639));
    InMux I__5454 (
            .O(N__29735),
            .I(N__29639));
    InMux I__5453 (
            .O(N__29734),
            .I(N__29639));
    InMux I__5452 (
            .O(N__29733),
            .I(N__29639));
    InMux I__5451 (
            .O(N__29732),
            .I(N__29634));
    InMux I__5450 (
            .O(N__29731),
            .I(N__29634));
    LocalMux I__5449 (
            .O(N__29722),
            .I(N__29631));
    LocalMux I__5448 (
            .O(N__29719),
            .I(N__29625));
    LocalMux I__5447 (
            .O(N__29710),
            .I(N__29625));
    InMux I__5446 (
            .O(N__29709),
            .I(N__29618));
    InMux I__5445 (
            .O(N__29708),
            .I(N__29618));
    InMux I__5444 (
            .O(N__29707),
            .I(N__29618));
    InMux I__5443 (
            .O(N__29706),
            .I(N__29609));
    InMux I__5442 (
            .O(N__29705),
            .I(N__29609));
    InMux I__5441 (
            .O(N__29704),
            .I(N__29609));
    InMux I__5440 (
            .O(N__29703),
            .I(N__29609));
    InMux I__5439 (
            .O(N__29702),
            .I(N__29600));
    InMux I__5438 (
            .O(N__29701),
            .I(N__29600));
    InMux I__5437 (
            .O(N__29700),
            .I(N__29600));
    InMux I__5436 (
            .O(N__29699),
            .I(N__29600));
    InMux I__5435 (
            .O(N__29698),
            .I(N__29595));
    InMux I__5434 (
            .O(N__29697),
            .I(N__29595));
    CascadeMux I__5433 (
            .O(N__29696),
            .I(N__29592));
    LocalMux I__5432 (
            .O(N__29693),
            .I(N__29588));
    InMux I__5431 (
            .O(N__29692),
            .I(N__29585));
    InMux I__5430 (
            .O(N__29691),
            .I(N__29582));
    InMux I__5429 (
            .O(N__29690),
            .I(N__29576));
    LocalMux I__5428 (
            .O(N__29687),
            .I(N__29573));
    LocalMux I__5427 (
            .O(N__29682),
            .I(N__29570));
    Span4Mux_v I__5426 (
            .O(N__29675),
            .I(N__29563));
    LocalMux I__5425 (
            .O(N__29670),
            .I(N__29563));
    Span4Mux_v I__5424 (
            .O(N__29665),
            .I(N__29563));
    LocalMux I__5423 (
            .O(N__29662),
            .I(N__29550));
    Span4Mux_v I__5422 (
            .O(N__29651),
            .I(N__29550));
    Span4Mux_h I__5421 (
            .O(N__29648),
            .I(N__29550));
    LocalMux I__5420 (
            .O(N__29639),
            .I(N__29550));
    LocalMux I__5419 (
            .O(N__29634),
            .I(N__29550));
    Span4Mux_h I__5418 (
            .O(N__29631),
            .I(N__29550));
    InMux I__5417 (
            .O(N__29630),
            .I(N__29547));
    Span4Mux_v I__5416 (
            .O(N__29625),
            .I(N__29536));
    LocalMux I__5415 (
            .O(N__29618),
            .I(N__29536));
    LocalMux I__5414 (
            .O(N__29609),
            .I(N__29536));
    LocalMux I__5413 (
            .O(N__29600),
            .I(N__29536));
    LocalMux I__5412 (
            .O(N__29595),
            .I(N__29536));
    InMux I__5411 (
            .O(N__29592),
            .I(N__29529));
    InMux I__5410 (
            .O(N__29591),
            .I(N__29529));
    Span4Mux_h I__5409 (
            .O(N__29588),
            .I(N__29524));
    LocalMux I__5408 (
            .O(N__29585),
            .I(N__29524));
    LocalMux I__5407 (
            .O(N__29582),
            .I(N__29521));
    InMux I__5406 (
            .O(N__29581),
            .I(N__29516));
    InMux I__5405 (
            .O(N__29580),
            .I(N__29516));
    InMux I__5404 (
            .O(N__29579),
            .I(N__29513));
    LocalMux I__5403 (
            .O(N__29576),
            .I(N__29504));
    Span4Mux_v I__5402 (
            .O(N__29573),
            .I(N__29504));
    Span4Mux_v I__5401 (
            .O(N__29570),
            .I(N__29504));
    Span4Mux_v I__5400 (
            .O(N__29563),
            .I(N__29504));
    Span4Mux_v I__5399 (
            .O(N__29550),
            .I(N__29501));
    LocalMux I__5398 (
            .O(N__29547),
            .I(N__29496));
    Span4Mux_v I__5397 (
            .O(N__29536),
            .I(N__29496));
    InMux I__5396 (
            .O(N__29535),
            .I(N__29491));
    InMux I__5395 (
            .O(N__29534),
            .I(N__29491));
    LocalMux I__5394 (
            .O(N__29529),
            .I(N__29484));
    Span4Mux_v I__5393 (
            .O(N__29524),
            .I(N__29484));
    Span4Mux_h I__5392 (
            .O(N__29521),
            .I(N__29484));
    LocalMux I__5391 (
            .O(N__29516),
            .I(N__29481));
    LocalMux I__5390 (
            .O(N__29513),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5389 (
            .O(N__29504),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5388 (
            .O(N__29501),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5387 (
            .O(N__29496),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__5386 (
            .O(N__29491),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5385 (
            .O(N__29484),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5384 (
            .O(N__29481),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__5383 (
            .O(N__29466),
            .I(N__29461));
    InMux I__5382 (
            .O(N__29465),
            .I(N__29458));
    InMux I__5381 (
            .O(N__29464),
            .I(N__29455));
    LocalMux I__5380 (
            .O(N__29461),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__5379 (
            .O(N__29458),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__5378 (
            .O(N__29455),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__5377 (
            .O(N__29448),
            .I(N__29445));
    LocalMux I__5376 (
            .O(N__29445),
            .I(N__29442));
    Span4Mux_h I__5375 (
            .O(N__29442),
            .I(N__29439));
    Span4Mux_v I__5374 (
            .O(N__29439),
            .I(N__29436));
    Odrv4 I__5373 (
            .O(N__29436),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__5372 (
            .O(N__29433),
            .I(N__29430));
    LocalMux I__5371 (
            .O(N__29430),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__5370 (
            .O(N__29427),
            .I(N__29424));
    LocalMux I__5369 (
            .O(N__29424),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__5368 (
            .O(N__29421),
            .I(N__29418));
    LocalMux I__5367 (
            .O(N__29418),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__5366 (
            .O(N__29415),
            .I(N__29412));
    LocalMux I__5365 (
            .O(N__29412),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__5364 (
            .O(N__29409),
            .I(N__29406));
    LocalMux I__5363 (
            .O(N__29406),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__5362 (
            .O(N__29403),
            .I(N__29400));
    LocalMux I__5361 (
            .O(N__29400),
            .I(N__29396));
    InMux I__5360 (
            .O(N__29399),
            .I(N__29393));
    Span4Mux_s1_v I__5359 (
            .O(N__29396),
            .I(N__29387));
    LocalMux I__5358 (
            .O(N__29393),
            .I(N__29387));
    InMux I__5357 (
            .O(N__29392),
            .I(N__29384));
    Span4Mux_v I__5356 (
            .O(N__29387),
            .I(N__29380));
    LocalMux I__5355 (
            .O(N__29384),
            .I(N__29377));
    InMux I__5354 (
            .O(N__29383),
            .I(N__29374));
    Span4Mux_h I__5353 (
            .O(N__29380),
            .I(N__29370));
    Span4Mux_h I__5352 (
            .O(N__29377),
            .I(N__29365));
    LocalMux I__5351 (
            .O(N__29374),
            .I(N__29365));
    InMux I__5350 (
            .O(N__29373),
            .I(N__29362));
    Sp12to4 I__5349 (
            .O(N__29370),
            .I(N__29359));
    Span4Mux_v I__5348 (
            .O(N__29365),
            .I(N__29356));
    LocalMux I__5347 (
            .O(N__29362),
            .I(N__29353));
    Span12Mux_v I__5346 (
            .O(N__29359),
            .I(N__29350));
    Sp12to4 I__5345 (
            .O(N__29356),
            .I(N__29347));
    Span4Mux_v I__5344 (
            .O(N__29353),
            .I(N__29344));
    Span12Mux_v I__5343 (
            .O(N__29350),
            .I(N__29341));
    Span12Mux_h I__5342 (
            .O(N__29347),
            .I(N__29338));
    Sp12to4 I__5341 (
            .O(N__29344),
            .I(N__29335));
    Span12Mux_h I__5340 (
            .O(N__29341),
            .I(N__29330));
    Span12Mux_v I__5339 (
            .O(N__29338),
            .I(N__29330));
    Span12Mux_h I__5338 (
            .O(N__29335),
            .I(N__29327));
    Odrv12 I__5337 (
            .O(N__29330),
            .I(start_stop_c));
    Odrv12 I__5336 (
            .O(N__29327),
            .I(start_stop_c));
    CEMux I__5335 (
            .O(N__29322),
            .I(N__29317));
    CEMux I__5334 (
            .O(N__29321),
            .I(N__29313));
    CEMux I__5333 (
            .O(N__29320),
            .I(N__29310));
    LocalMux I__5332 (
            .O(N__29317),
            .I(N__29307));
    CEMux I__5331 (
            .O(N__29316),
            .I(N__29304));
    LocalMux I__5330 (
            .O(N__29313),
            .I(N__29301));
    LocalMux I__5329 (
            .O(N__29310),
            .I(N__29298));
    Span4Mux_h I__5328 (
            .O(N__29307),
            .I(N__29295));
    LocalMux I__5327 (
            .O(N__29304),
            .I(N__29292));
    Span4Mux_h I__5326 (
            .O(N__29301),
            .I(N__29289));
    Span4Mux_v I__5325 (
            .O(N__29298),
            .I(N__29286));
    Span4Mux_v I__5324 (
            .O(N__29295),
            .I(N__29281));
    Span4Mux_h I__5323 (
            .O(N__29292),
            .I(N__29281));
    Sp12to4 I__5322 (
            .O(N__29289),
            .I(N__29277));
    Span4Mux_v I__5321 (
            .O(N__29286),
            .I(N__29274));
    Span4Mux_v I__5320 (
            .O(N__29281),
            .I(N__29271));
    CEMux I__5319 (
            .O(N__29280),
            .I(N__29268));
    Odrv12 I__5318 (
            .O(N__29277),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__5317 (
            .O(N__29274),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    Odrv4 I__5316 (
            .O(N__29271),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    LocalMux I__5315 (
            .O(N__29268),
            .I(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ));
    InMux I__5314 (
            .O(N__29259),
            .I(N__29256));
    LocalMux I__5313 (
            .O(N__29256),
            .I(N__29253));
    Span4Mux_v I__5312 (
            .O(N__29253),
            .I(N__29248));
    InMux I__5311 (
            .O(N__29252),
            .I(N__29245));
    InMux I__5310 (
            .O(N__29251),
            .I(N__29242));
    Odrv4 I__5309 (
            .O(N__29248),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__5308 (
            .O(N__29245),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__5307 (
            .O(N__29242),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__5306 (
            .O(N__29235),
            .I(N__29232));
    LocalMux I__5305 (
            .O(N__29232),
            .I(N__29229));
    Span4Mux_v I__5304 (
            .O(N__29229),
            .I(N__29226));
    Span4Mux_h I__5303 (
            .O(N__29226),
            .I(N__29223));
    Odrv4 I__5302 (
            .O(N__29223),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__5301 (
            .O(N__29220),
            .I(N__29217));
    LocalMux I__5300 (
            .O(N__29217),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__5299 (
            .O(N__29214),
            .I(N__29208));
    InMux I__5298 (
            .O(N__29213),
            .I(N__29205));
    InMux I__5297 (
            .O(N__29212),
            .I(N__29200));
    InMux I__5296 (
            .O(N__29211),
            .I(N__29200));
    LocalMux I__5295 (
            .O(N__29208),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__5294 (
            .O(N__29205),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__5293 (
            .O(N__29200),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__5292 (
            .O(N__29193),
            .I(N__29190));
    LocalMux I__5291 (
            .O(N__29190),
            .I(N__29186));
    InMux I__5290 (
            .O(N__29189),
            .I(N__29183));
    Span4Mux_h I__5289 (
            .O(N__29186),
            .I(N__29176));
    LocalMux I__5288 (
            .O(N__29183),
            .I(N__29176));
    InMux I__5287 (
            .O(N__29182),
            .I(N__29171));
    InMux I__5286 (
            .O(N__29181),
            .I(N__29171));
    Span4Mux_h I__5285 (
            .O(N__29176),
            .I(N__29168));
    LocalMux I__5284 (
            .O(N__29171),
            .I(N__29165));
    Odrv4 I__5283 (
            .O(N__29168),
            .I(\phase_controller_inst2.stoper_tr.time_passed11 ));
    Odrv12 I__5282 (
            .O(N__29165),
            .I(\phase_controller_inst2.stoper_tr.time_passed11 ));
    InMux I__5281 (
            .O(N__29160),
            .I(N__29153));
    InMux I__5280 (
            .O(N__29159),
            .I(N__29153));
    InMux I__5279 (
            .O(N__29158),
            .I(N__29149));
    LocalMux I__5278 (
            .O(N__29153),
            .I(N__29144));
    InMux I__5277 (
            .O(N__29152),
            .I(N__29141));
    LocalMux I__5276 (
            .O(N__29149),
            .I(N__29138));
    InMux I__5275 (
            .O(N__29148),
            .I(N__29133));
    InMux I__5274 (
            .O(N__29147),
            .I(N__29133));
    Span4Mux_h I__5273 (
            .O(N__29144),
            .I(N__29130));
    LocalMux I__5272 (
            .O(N__29141),
            .I(N__29127));
    Span4Mux_v I__5271 (
            .O(N__29138),
            .I(N__29122));
    LocalMux I__5270 (
            .O(N__29133),
            .I(N__29122));
    Odrv4 I__5269 (
            .O(N__29130),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__5268 (
            .O(N__29127),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    Odrv4 I__5267 (
            .O(N__29122),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ));
    CascadeMux I__5266 (
            .O(N__29115),
            .I(N__29112));
    InMux I__5265 (
            .O(N__29112),
            .I(N__29105));
    InMux I__5264 (
            .O(N__29111),
            .I(N__29105));
    CascadeMux I__5263 (
            .O(N__29110),
            .I(N__29095));
    LocalMux I__5262 (
            .O(N__29105),
            .I(N__29091));
    InMux I__5261 (
            .O(N__29104),
            .I(N__29088));
    InMux I__5260 (
            .O(N__29103),
            .I(N__29068));
    InMux I__5259 (
            .O(N__29102),
            .I(N__29068));
    InMux I__5258 (
            .O(N__29101),
            .I(N__29068));
    InMux I__5257 (
            .O(N__29100),
            .I(N__29068));
    InMux I__5256 (
            .O(N__29099),
            .I(N__29068));
    InMux I__5255 (
            .O(N__29098),
            .I(N__29068));
    InMux I__5254 (
            .O(N__29095),
            .I(N__29068));
    InMux I__5253 (
            .O(N__29094),
            .I(N__29065));
    Span4Mux_v I__5252 (
            .O(N__29091),
            .I(N__29060));
    LocalMux I__5251 (
            .O(N__29088),
            .I(N__29060));
    CascadeMux I__5250 (
            .O(N__29087),
            .I(N__29055));
    CascadeMux I__5249 (
            .O(N__29086),
            .I(N__29052));
    CascadeMux I__5248 (
            .O(N__29085),
            .I(N__29049));
    CascadeMux I__5247 (
            .O(N__29084),
            .I(N__29043));
    CascadeMux I__5246 (
            .O(N__29083),
            .I(N__29040));
    LocalMux I__5245 (
            .O(N__29068),
            .I(N__29034));
    LocalMux I__5244 (
            .O(N__29065),
            .I(N__29029));
    Span4Mux_h I__5243 (
            .O(N__29060),
            .I(N__29029));
    InMux I__5242 (
            .O(N__29059),
            .I(N__29026));
    InMux I__5241 (
            .O(N__29058),
            .I(N__29023));
    InMux I__5240 (
            .O(N__29055),
            .I(N__29010));
    InMux I__5239 (
            .O(N__29052),
            .I(N__29010));
    InMux I__5238 (
            .O(N__29049),
            .I(N__29010));
    InMux I__5237 (
            .O(N__29048),
            .I(N__29010));
    InMux I__5236 (
            .O(N__29047),
            .I(N__29010));
    InMux I__5235 (
            .O(N__29046),
            .I(N__29010));
    InMux I__5234 (
            .O(N__29043),
            .I(N__29003));
    InMux I__5233 (
            .O(N__29040),
            .I(N__29003));
    InMux I__5232 (
            .O(N__29039),
            .I(N__29003));
    InMux I__5231 (
            .O(N__29038),
            .I(N__28998));
    InMux I__5230 (
            .O(N__29037),
            .I(N__28998));
    Span4Mux_h I__5229 (
            .O(N__29034),
            .I(N__28993));
    Span4Mux_h I__5228 (
            .O(N__29029),
            .I(N__28993));
    LocalMux I__5227 (
            .O(N__29026),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__5226 (
            .O(N__29023),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__5225 (
            .O(N__29010),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__5224 (
            .O(N__29003),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__5223 (
            .O(N__28998),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__5222 (
            .O(N__28993),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CascadeMux I__5221 (
            .O(N__28980),
            .I(N__28975));
    CascadeMux I__5220 (
            .O(N__28979),
            .I(N__28972));
    CascadeMux I__5219 (
            .O(N__28978),
            .I(N__28969));
    InMux I__5218 (
            .O(N__28975),
            .I(N__28956));
    InMux I__5217 (
            .O(N__28972),
            .I(N__28956));
    InMux I__5216 (
            .O(N__28969),
            .I(N__28956));
    CascadeMux I__5215 (
            .O(N__28968),
            .I(N__28953));
    CascadeMux I__5214 (
            .O(N__28967),
            .I(N__28950));
    CascadeMux I__5213 (
            .O(N__28966),
            .I(N__28947));
    CascadeMux I__5212 (
            .O(N__28965),
            .I(N__28938));
    InMux I__5211 (
            .O(N__28964),
            .I(N__28928));
    InMux I__5210 (
            .O(N__28963),
            .I(N__28928));
    LocalMux I__5209 (
            .O(N__28956),
            .I(N__28924));
    InMux I__5208 (
            .O(N__28953),
            .I(N__28913));
    InMux I__5207 (
            .O(N__28950),
            .I(N__28913));
    InMux I__5206 (
            .O(N__28947),
            .I(N__28913));
    InMux I__5205 (
            .O(N__28946),
            .I(N__28913));
    InMux I__5204 (
            .O(N__28945),
            .I(N__28913));
    InMux I__5203 (
            .O(N__28944),
            .I(N__28906));
    InMux I__5202 (
            .O(N__28943),
            .I(N__28906));
    InMux I__5201 (
            .O(N__28942),
            .I(N__28906));
    InMux I__5200 (
            .O(N__28941),
            .I(N__28891));
    InMux I__5199 (
            .O(N__28938),
            .I(N__28891));
    InMux I__5198 (
            .O(N__28937),
            .I(N__28891));
    InMux I__5197 (
            .O(N__28936),
            .I(N__28891));
    InMux I__5196 (
            .O(N__28935),
            .I(N__28891));
    InMux I__5195 (
            .O(N__28934),
            .I(N__28891));
    InMux I__5194 (
            .O(N__28933),
            .I(N__28891));
    LocalMux I__5193 (
            .O(N__28928),
            .I(N__28888));
    CascadeMux I__5192 (
            .O(N__28927),
            .I(N__28884));
    Span4Mux_v I__5191 (
            .O(N__28924),
            .I(N__28878));
    LocalMux I__5190 (
            .O(N__28913),
            .I(N__28878));
    LocalMux I__5189 (
            .O(N__28906),
            .I(N__28875));
    LocalMux I__5188 (
            .O(N__28891),
            .I(N__28870));
    Span4Mux_h I__5187 (
            .O(N__28888),
            .I(N__28870));
    InMux I__5186 (
            .O(N__28887),
            .I(N__28867));
    InMux I__5185 (
            .O(N__28884),
            .I(N__28861));
    InMux I__5184 (
            .O(N__28883),
            .I(N__28861));
    Span4Mux_h I__5183 (
            .O(N__28878),
            .I(N__28858));
    Span4Mux_h I__5182 (
            .O(N__28875),
            .I(N__28855));
    Span4Mux_h I__5181 (
            .O(N__28870),
            .I(N__28850));
    LocalMux I__5180 (
            .O(N__28867),
            .I(N__28850));
    InMux I__5179 (
            .O(N__28866),
            .I(N__28847));
    LocalMux I__5178 (
            .O(N__28861),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__5177 (
            .O(N__28858),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__5176 (
            .O(N__28855),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    Odrv4 I__5175 (
            .O(N__28850),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    LocalMux I__5174 (
            .O(N__28847),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ));
    CascadeMux I__5173 (
            .O(N__28836),
            .I(N__28833));
    InMux I__5172 (
            .O(N__28833),
            .I(N__28797));
    InMux I__5171 (
            .O(N__28832),
            .I(N__28797));
    InMux I__5170 (
            .O(N__28831),
            .I(N__28797));
    InMux I__5169 (
            .O(N__28830),
            .I(N__28797));
    InMux I__5168 (
            .O(N__28829),
            .I(N__28797));
    InMux I__5167 (
            .O(N__28828),
            .I(N__28797));
    InMux I__5166 (
            .O(N__28827),
            .I(N__28797));
    InMux I__5165 (
            .O(N__28826),
            .I(N__28797));
    InMux I__5164 (
            .O(N__28825),
            .I(N__28790));
    InMux I__5163 (
            .O(N__28824),
            .I(N__28790));
    InMux I__5162 (
            .O(N__28823),
            .I(N__28790));
    InMux I__5161 (
            .O(N__28822),
            .I(N__28785));
    InMux I__5160 (
            .O(N__28821),
            .I(N__28785));
    InMux I__5159 (
            .O(N__28820),
            .I(N__28770));
    InMux I__5158 (
            .O(N__28819),
            .I(N__28770));
    InMux I__5157 (
            .O(N__28818),
            .I(N__28770));
    InMux I__5156 (
            .O(N__28817),
            .I(N__28770));
    InMux I__5155 (
            .O(N__28816),
            .I(N__28770));
    InMux I__5154 (
            .O(N__28815),
            .I(N__28770));
    InMux I__5153 (
            .O(N__28814),
            .I(N__28770));
    LocalMux I__5152 (
            .O(N__28797),
            .I(N__28764));
    LocalMux I__5151 (
            .O(N__28790),
            .I(N__28761));
    LocalMux I__5150 (
            .O(N__28785),
            .I(N__28758));
    LocalMux I__5149 (
            .O(N__28770),
            .I(N__28755));
    InMux I__5148 (
            .O(N__28769),
            .I(N__28752));
    InMux I__5147 (
            .O(N__28768),
            .I(N__28746));
    InMux I__5146 (
            .O(N__28767),
            .I(N__28746));
    Span4Mux_h I__5145 (
            .O(N__28764),
            .I(N__28743));
    Span4Mux_h I__5144 (
            .O(N__28761),
            .I(N__28740));
    Span12Mux_v I__5143 (
            .O(N__28758),
            .I(N__28737));
    Span4Mux_h I__5142 (
            .O(N__28755),
            .I(N__28732));
    LocalMux I__5141 (
            .O(N__28752),
            .I(N__28732));
    InMux I__5140 (
            .O(N__28751),
            .I(N__28729));
    LocalMux I__5139 (
            .O(N__28746),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__5138 (
            .O(N__28743),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__5137 (
            .O(N__28740),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv12 I__5136 (
            .O(N__28737),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    Odrv4 I__5135 (
            .O(N__28732),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    LocalMux I__5134 (
            .O(N__28729),
            .I(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ));
    InMux I__5133 (
            .O(N__28716),
            .I(N__28713));
    LocalMux I__5132 (
            .O(N__28713),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__5131 (
            .O(N__28710),
            .I(N__28707));
    LocalMux I__5130 (
            .O(N__28707),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__5129 (
            .O(N__28704),
            .I(N__28700));
    CascadeMux I__5128 (
            .O(N__28703),
            .I(N__28695));
    LocalMux I__5127 (
            .O(N__28700),
            .I(N__28688));
    InMux I__5126 (
            .O(N__28699),
            .I(N__28677));
    InMux I__5125 (
            .O(N__28698),
            .I(N__28677));
    InMux I__5124 (
            .O(N__28695),
            .I(N__28677));
    InMux I__5123 (
            .O(N__28694),
            .I(N__28677));
    InMux I__5122 (
            .O(N__28693),
            .I(N__28672));
    InMux I__5121 (
            .O(N__28692),
            .I(N__28672));
    CascadeMux I__5120 (
            .O(N__28691),
            .I(N__28668));
    Span4Mux_h I__5119 (
            .O(N__28688),
            .I(N__28664));
    InMux I__5118 (
            .O(N__28687),
            .I(N__28659));
    InMux I__5117 (
            .O(N__28686),
            .I(N__28659));
    LocalMux I__5116 (
            .O(N__28677),
            .I(N__28654));
    LocalMux I__5115 (
            .O(N__28672),
            .I(N__28654));
    InMux I__5114 (
            .O(N__28671),
            .I(N__28647));
    InMux I__5113 (
            .O(N__28668),
            .I(N__28647));
    InMux I__5112 (
            .O(N__28667),
            .I(N__28647));
    Odrv4 I__5111 (
            .O(N__28664),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__5110 (
            .O(N__28659),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    Odrv4 I__5109 (
            .O(N__28654),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    LocalMux I__5108 (
            .O(N__28647),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ));
    InMux I__5107 (
            .O(N__28638),
            .I(N__28635));
    LocalMux I__5106 (
            .O(N__28635),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ));
    InMux I__5105 (
            .O(N__28632),
            .I(N__28629));
    LocalMux I__5104 (
            .O(N__28629),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ));
    CascadeMux I__5103 (
            .O(N__28626),
            .I(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ));
    InMux I__5102 (
            .O(N__28623),
            .I(N__28620));
    LocalMux I__5101 (
            .O(N__28620),
            .I(N__28616));
    InMux I__5100 (
            .O(N__28619),
            .I(N__28613));
    Odrv4 I__5099 (
            .O(N__28616),
            .I(\phase_controller_inst1.stoper_tr.N_257 ));
    LocalMux I__5098 (
            .O(N__28613),
            .I(\phase_controller_inst1.stoper_tr.N_257 ));
    CascadeMux I__5097 (
            .O(N__28608),
            .I(\phase_controller_inst1.stoper_tr.N_257_cascade_ ));
    InMux I__5096 (
            .O(N__28605),
            .I(N__28599));
    InMux I__5095 (
            .O(N__28604),
            .I(N__28599));
    LocalMux I__5094 (
            .O(N__28599),
            .I(N__28594));
    InMux I__5093 (
            .O(N__28598),
            .I(N__28589));
    InMux I__5092 (
            .O(N__28597),
            .I(N__28589));
    Odrv4 I__5091 (
            .O(N__28594),
            .I(\phase_controller_inst1.stoper_tr.N_240 ));
    LocalMux I__5090 (
            .O(N__28589),
            .I(\phase_controller_inst1.stoper_tr.N_240 ));
    InMux I__5089 (
            .O(N__28584),
            .I(N__28578));
    InMux I__5088 (
            .O(N__28583),
            .I(N__28578));
    LocalMux I__5087 (
            .O(N__28578),
            .I(N__28574));
    InMux I__5086 (
            .O(N__28577),
            .I(N__28571));
    Odrv12 I__5085 (
            .O(N__28574),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__5084 (
            .O(N__28571),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__5083 (
            .O(N__28566),
            .I(N__28563));
    LocalMux I__5082 (
            .O(N__28563),
            .I(N__28560));
    Odrv4 I__5081 (
            .O(N__28560),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__5080 (
            .O(N__28557),
            .I(N__28554));
    LocalMux I__5079 (
            .O(N__28554),
            .I(N__28551));
    Span4Mux_v I__5078 (
            .O(N__28551),
            .I(N__28548));
    Odrv4 I__5077 (
            .O(N__28548),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__5076 (
            .O(N__28545),
            .I(N__28541));
    InMux I__5075 (
            .O(N__28544),
            .I(N__28538));
    LocalMux I__5074 (
            .O(N__28541),
            .I(N__28535));
    LocalMux I__5073 (
            .O(N__28538),
            .I(N__28532));
    Odrv4 I__5072 (
            .O(N__28535),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    Odrv12 I__5071 (
            .O(N__28532),
            .I(\current_shift_inst.un4_control_input_0_31 ));
    IoInMux I__5070 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__5069 (
            .O(N__28524),
            .I(N__28521));
    Odrv12 I__5068 (
            .O(N__28521),
            .I(\delay_measurement_inst.delay_tr_timer.N_463_i ));
    InMux I__5067 (
            .O(N__28518),
            .I(N__28514));
    InMux I__5066 (
            .O(N__28517),
            .I(N__28511));
    LocalMux I__5065 (
            .O(N__28514),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__5064 (
            .O(N__28511),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__5063 (
            .O(N__28506),
            .I(N__28502));
    InMux I__5062 (
            .O(N__28505),
            .I(N__28498));
    LocalMux I__5061 (
            .O(N__28502),
            .I(N__28495));
    InMux I__5060 (
            .O(N__28501),
            .I(N__28492));
    LocalMux I__5059 (
            .O(N__28498),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__5058 (
            .O(N__28495),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__5057 (
            .O(N__28492),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__5056 (
            .O(N__28485),
            .I(N__28482));
    LocalMux I__5055 (
            .O(N__28482),
            .I(N__28478));
    InMux I__5054 (
            .O(N__28481),
            .I(N__28475));
    Sp12to4 I__5053 (
            .O(N__28478),
            .I(N__28469));
    LocalMux I__5052 (
            .O(N__28475),
            .I(N__28469));
    InMux I__5051 (
            .O(N__28474),
            .I(N__28466));
    Odrv12 I__5050 (
            .O(N__28469),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__5049 (
            .O(N__28466),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__5048 (
            .O(N__28461),
            .I(N__28458));
    LocalMux I__5047 (
            .O(N__28458),
            .I(N__28455));
    Span4Mux_h I__5046 (
            .O(N__28455),
            .I(N__28452));
    Odrv4 I__5045 (
            .O(N__28452),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__5044 (
            .O(N__28449),
            .I(N__28446));
    LocalMux I__5043 (
            .O(N__28446),
            .I(N__28443));
    Span4Mux_v I__5042 (
            .O(N__28443),
            .I(N__28440));
    Odrv4 I__5041 (
            .O(N__28440),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__5040 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__5039 (
            .O(N__28434),
            .I(N__28430));
    InMux I__5038 (
            .O(N__28433),
            .I(N__28427));
    Sp12to4 I__5037 (
            .O(N__28430),
            .I(N__28421));
    LocalMux I__5036 (
            .O(N__28427),
            .I(N__28421));
    InMux I__5035 (
            .O(N__28426),
            .I(N__28418));
    Odrv12 I__5034 (
            .O(N__28421),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__5033 (
            .O(N__28418),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__5032 (
            .O(N__28413),
            .I(N__28410));
    LocalMux I__5031 (
            .O(N__28410),
            .I(N__28407));
    Odrv4 I__5030 (
            .O(N__28407),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__5029 (
            .O(N__28404),
            .I(N__28401));
    LocalMux I__5028 (
            .O(N__28401),
            .I(N__28396));
    InMux I__5027 (
            .O(N__28400),
            .I(N__28391));
    InMux I__5026 (
            .O(N__28399),
            .I(N__28391));
    Odrv4 I__5025 (
            .O(N__28396),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__5024 (
            .O(N__28391),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__5023 (
            .O(N__28386),
            .I(N__28383));
    LocalMux I__5022 (
            .O(N__28383),
            .I(N__28380));
    Span4Mux_h I__5021 (
            .O(N__28380),
            .I(N__28377));
    Odrv4 I__5020 (
            .O(N__28377),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__5019 (
            .O(N__28374),
            .I(N__28371));
    LocalMux I__5018 (
            .O(N__28371),
            .I(N__28367));
    InMux I__5017 (
            .O(N__28370),
            .I(N__28364));
    Sp12to4 I__5016 (
            .O(N__28367),
            .I(N__28358));
    LocalMux I__5015 (
            .O(N__28364),
            .I(N__28358));
    InMux I__5014 (
            .O(N__28363),
            .I(N__28355));
    Odrv12 I__5013 (
            .O(N__28358),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__5012 (
            .O(N__28355),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__5011 (
            .O(N__28350),
            .I(N__28347));
    LocalMux I__5010 (
            .O(N__28347),
            .I(N__28344));
    Odrv12 I__5009 (
            .O(N__28344),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__5008 (
            .O(N__28341),
            .I(N__28338));
    LocalMux I__5007 (
            .O(N__28338),
            .I(N__28334));
    InMux I__5006 (
            .O(N__28337),
            .I(N__28331));
    Sp12to4 I__5005 (
            .O(N__28334),
            .I(N__28325));
    LocalMux I__5004 (
            .O(N__28331),
            .I(N__28325));
    InMux I__5003 (
            .O(N__28330),
            .I(N__28322));
    Odrv12 I__5002 (
            .O(N__28325),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__5001 (
            .O(N__28322),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__5000 (
            .O(N__28317),
            .I(N__28314));
    LocalMux I__4999 (
            .O(N__28314),
            .I(N__28311));
    Odrv4 I__4998 (
            .O(N__28311),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__4997 (
            .O(N__28308),
            .I(N__28305));
    LocalMux I__4996 (
            .O(N__28305),
            .I(N__28301));
    InMux I__4995 (
            .O(N__28304),
            .I(N__28298));
    Span4Mux_v I__4994 (
            .O(N__28301),
            .I(N__28294));
    LocalMux I__4993 (
            .O(N__28298),
            .I(N__28291));
    InMux I__4992 (
            .O(N__28297),
            .I(N__28288));
    Odrv4 I__4991 (
            .O(N__28294),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv12 I__4990 (
            .O(N__28291),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__4989 (
            .O(N__28288),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__4988 (
            .O(N__28281),
            .I(N__28278));
    LocalMux I__4987 (
            .O(N__28278),
            .I(N__28275));
    Odrv4 I__4986 (
            .O(N__28275),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__4985 (
            .O(N__28272),
            .I(N__28269));
    LocalMux I__4984 (
            .O(N__28269),
            .I(N__28265));
    InMux I__4983 (
            .O(N__28268),
            .I(N__28262));
    Span4Mux_v I__4982 (
            .O(N__28265),
            .I(N__28258));
    LocalMux I__4981 (
            .O(N__28262),
            .I(N__28255));
    InMux I__4980 (
            .O(N__28261),
            .I(N__28252));
    Odrv4 I__4979 (
            .O(N__28258),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv12 I__4978 (
            .O(N__28255),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__4977 (
            .O(N__28252),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__4976 (
            .O(N__28245),
            .I(N__28242));
    LocalMux I__4975 (
            .O(N__28242),
            .I(N__28239));
    Odrv4 I__4974 (
            .O(N__28239),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__4973 (
            .O(N__28236),
            .I(N__28233));
    LocalMux I__4972 (
            .O(N__28233),
            .I(N__28230));
    Odrv4 I__4971 (
            .O(N__28230),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    CascadeMux I__4970 (
            .O(N__28227),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__4969 (
            .O(N__28224),
            .I(N__28221));
    LocalMux I__4968 (
            .O(N__28221),
            .I(N__28218));
    Span4Mux_h I__4967 (
            .O(N__28218),
            .I(N__28215));
    Odrv4 I__4966 (
            .O(N__28215),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__4965 (
            .O(N__28212),
            .I(N__28209));
    LocalMux I__4964 (
            .O(N__28209),
            .I(N__28206));
    Span4Mux_v I__4963 (
            .O(N__28206),
            .I(N__28201));
    InMux I__4962 (
            .O(N__28205),
            .I(N__28198));
    InMux I__4961 (
            .O(N__28204),
            .I(N__28195));
    Odrv4 I__4960 (
            .O(N__28201),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__4959 (
            .O(N__28198),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__4958 (
            .O(N__28195),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__4957 (
            .O(N__28188),
            .I(N__28185));
    LocalMux I__4956 (
            .O(N__28185),
            .I(N__28182));
    Span12Mux_v I__4955 (
            .O(N__28182),
            .I(N__28179));
    Odrv12 I__4954 (
            .O(N__28179),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__4953 (
            .O(N__28176),
            .I(N__28173));
    LocalMux I__4952 (
            .O(N__28173),
            .I(N__28170));
    Span4Mux_v I__4951 (
            .O(N__28170),
            .I(N__28167));
    Odrv4 I__4950 (
            .O(N__28167),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__4949 (
            .O(N__28164),
            .I(N__28161));
    LocalMux I__4948 (
            .O(N__28161),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__4947 (
            .O(N__28158),
            .I(N__28155));
    LocalMux I__4946 (
            .O(N__28155),
            .I(N__28152));
    Span4Mux_h I__4945 (
            .O(N__28152),
            .I(N__28149));
    Span4Mux_v I__4944 (
            .O(N__28149),
            .I(N__28146));
    Odrv4 I__4943 (
            .O(N__28146),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__4942 (
            .O(N__28143),
            .I(N__28134));
    InMux I__4941 (
            .O(N__28142),
            .I(N__28134));
    InMux I__4940 (
            .O(N__28141),
            .I(N__28134));
    LocalMux I__4939 (
            .O(N__28134),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__4938 (
            .O(N__28131),
            .I(N__28128));
    LocalMux I__4937 (
            .O(N__28128),
            .I(N__28125));
    Odrv4 I__4936 (
            .O(N__28125),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__4935 (
            .O(N__28122),
            .I(N__28119));
    LocalMux I__4934 (
            .O(N__28119),
            .I(N__28115));
    InMux I__4933 (
            .O(N__28118),
            .I(N__28112));
    Span4Mux_v I__4932 (
            .O(N__28115),
            .I(N__28106));
    LocalMux I__4931 (
            .O(N__28112),
            .I(N__28106));
    InMux I__4930 (
            .O(N__28111),
            .I(N__28103));
    Odrv4 I__4929 (
            .O(N__28106),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__4928 (
            .O(N__28103),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__4927 (
            .O(N__28098),
            .I(N__28095));
    LocalMux I__4926 (
            .O(N__28095),
            .I(N__28092));
    Span4Mux_h I__4925 (
            .O(N__28092),
            .I(N__28089));
    Odrv4 I__4924 (
            .O(N__28089),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__4923 (
            .O(N__28086),
            .I(N__28083));
    LocalMux I__4922 (
            .O(N__28083),
            .I(N__28079));
    InMux I__4921 (
            .O(N__28082),
            .I(N__28076));
    Span4Mux_v I__4920 (
            .O(N__28079),
            .I(N__28070));
    LocalMux I__4919 (
            .O(N__28076),
            .I(N__28070));
    InMux I__4918 (
            .O(N__28075),
            .I(N__28067));
    Odrv4 I__4917 (
            .O(N__28070),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__4916 (
            .O(N__28067),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__4915 (
            .O(N__28062),
            .I(N__28059));
    LocalMux I__4914 (
            .O(N__28059),
            .I(N__28056));
    Span4Mux_h I__4913 (
            .O(N__28056),
            .I(N__28053));
    Odrv4 I__4912 (
            .O(N__28053),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__4911 (
            .O(N__28050),
            .I(N__28047));
    LocalMux I__4910 (
            .O(N__28047),
            .I(N__28043));
    InMux I__4909 (
            .O(N__28046),
            .I(N__28040));
    Span4Mux_v I__4908 (
            .O(N__28043),
            .I(N__28034));
    LocalMux I__4907 (
            .O(N__28040),
            .I(N__28034));
    InMux I__4906 (
            .O(N__28039),
            .I(N__28031));
    Odrv4 I__4905 (
            .O(N__28034),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__4904 (
            .O(N__28031),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__4903 (
            .O(N__28026),
            .I(N__28023));
    LocalMux I__4902 (
            .O(N__28023),
            .I(N__28020));
    Span4Mux_h I__4901 (
            .O(N__28020),
            .I(N__28017));
    Odrv4 I__4900 (
            .O(N__28017),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__4899 (
            .O(N__28014),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__4898 (
            .O(N__28011),
            .I(N__28008));
    LocalMux I__4897 (
            .O(N__28008),
            .I(N__28005));
    Odrv12 I__4896 (
            .O(N__28005),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__4895 (
            .O(N__28002),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__4894 (
            .O(N__27999),
            .I(N__27992));
    InMux I__4893 (
            .O(N__27998),
            .I(N__27992));
    InMux I__4892 (
            .O(N__27997),
            .I(N__27989));
    LocalMux I__4891 (
            .O(N__27992),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__4890 (
            .O(N__27989),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__4889 (
            .O(N__27984),
            .I(bfn_11_17_0_));
    InMux I__4888 (
            .O(N__27981),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__4887 (
            .O(N__27978),
            .I(N__27975));
    LocalMux I__4886 (
            .O(N__27975),
            .I(N__27970));
    InMux I__4885 (
            .O(N__27974),
            .I(N__27965));
    InMux I__4884 (
            .O(N__27973),
            .I(N__27965));
    Odrv4 I__4883 (
            .O(N__27970),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__4882 (
            .O(N__27965),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__4881 (
            .O(N__27960),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__4880 (
            .O(N__27957),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__4879 (
            .O(N__27954),
            .I(N__27951));
    LocalMux I__4878 (
            .O(N__27951),
            .I(N__27947));
    InMux I__4877 (
            .O(N__27950),
            .I(N__27944));
    Span4Mux_v I__4876 (
            .O(N__27947),
            .I(N__27938));
    LocalMux I__4875 (
            .O(N__27944),
            .I(N__27938));
    InMux I__4874 (
            .O(N__27943),
            .I(N__27935));
    Odrv4 I__4873 (
            .O(N__27938),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__4872 (
            .O(N__27935),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__4871 (
            .O(N__27930),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__4870 (
            .O(N__27927),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__4869 (
            .O(N__27924),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__4868 (
            .O(N__27921),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__4867 (
            .O(N__27918),
            .I(N__27915));
    LocalMux I__4866 (
            .O(N__27915),
            .I(N__27912));
    Odrv4 I__4865 (
            .O(N__27912),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__4864 (
            .O(N__27909),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__4863 (
            .O(N__27906),
            .I(N__27903));
    LocalMux I__4862 (
            .O(N__27903),
            .I(N__27900));
    Odrv4 I__4861 (
            .O(N__27900),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__4860 (
            .O(N__27897),
            .I(N__27894));
    LocalMux I__4859 (
            .O(N__27894),
            .I(N__27890));
    InMux I__4858 (
            .O(N__27893),
            .I(N__27887));
    Span4Mux_h I__4857 (
            .O(N__27890),
            .I(N__27882));
    LocalMux I__4856 (
            .O(N__27887),
            .I(N__27882));
    Span4Mux_v I__4855 (
            .O(N__27882),
            .I(N__27878));
    InMux I__4854 (
            .O(N__27881),
            .I(N__27875));
    Odrv4 I__4853 (
            .O(N__27878),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__4852 (
            .O(N__27875),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__4851 (
            .O(N__27870),
            .I(bfn_11_16_0_));
    InMux I__4850 (
            .O(N__27867),
            .I(N__27864));
    LocalMux I__4849 (
            .O(N__27864),
            .I(N__27859));
    InMux I__4848 (
            .O(N__27863),
            .I(N__27854));
    InMux I__4847 (
            .O(N__27862),
            .I(N__27854));
    Odrv12 I__4846 (
            .O(N__27859),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__4845 (
            .O(N__27854),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__4844 (
            .O(N__27849),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__4843 (
            .O(N__27846),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__4842 (
            .O(N__27843),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__4841 (
            .O(N__27840),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__4840 (
            .O(N__27837),
            .I(N__27831));
    InMux I__4839 (
            .O(N__27836),
            .I(N__27831));
    LocalMux I__4838 (
            .O(N__27831),
            .I(N__27828));
    Span4Mux_v I__4837 (
            .O(N__27828),
            .I(N__27824));
    InMux I__4836 (
            .O(N__27827),
            .I(N__27821));
    Odrv4 I__4835 (
            .O(N__27824),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__4834 (
            .O(N__27821),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__4833 (
            .O(N__27816),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__4832 (
            .O(N__27813),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__4831 (
            .O(N__27810),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__4830 (
            .O(N__27807),
            .I(N__27803));
    InMux I__4829 (
            .O(N__27806),
            .I(N__27800));
    LocalMux I__4828 (
            .O(N__27803),
            .I(N__27797));
    LocalMux I__4827 (
            .O(N__27800),
            .I(N__27794));
    Span4Mux_v I__4826 (
            .O(N__27797),
            .I(N__27790));
    Span4Mux_v I__4825 (
            .O(N__27794),
            .I(N__27787));
    InMux I__4824 (
            .O(N__27793),
            .I(N__27784));
    Odrv4 I__4823 (
            .O(N__27790),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__4822 (
            .O(N__27787),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__4821 (
            .O(N__27784),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__4820 (
            .O(N__27777),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__4819 (
            .O(N__27774),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__4818 (
            .O(N__27771),
            .I(N__27768));
    LocalMux I__4817 (
            .O(N__27768),
            .I(N__27765));
    Span4Mux_h I__4816 (
            .O(N__27765),
            .I(N__27760));
    InMux I__4815 (
            .O(N__27764),
            .I(N__27757));
    InMux I__4814 (
            .O(N__27763),
            .I(N__27754));
    Odrv4 I__4813 (
            .O(N__27760),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__4812 (
            .O(N__27757),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__4811 (
            .O(N__27754),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__4810 (
            .O(N__27747),
            .I(bfn_11_15_0_));
    InMux I__4809 (
            .O(N__27744),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__4808 (
            .O(N__27741),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__4807 (
            .O(N__27738),
            .I(N__27735));
    LocalMux I__4806 (
            .O(N__27735),
            .I(N__27732));
    Span4Mux_v I__4805 (
            .O(N__27732),
            .I(N__27727));
    InMux I__4804 (
            .O(N__27731),
            .I(N__27724));
    InMux I__4803 (
            .O(N__27730),
            .I(N__27721));
    Odrv4 I__4802 (
            .O(N__27727),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__4801 (
            .O(N__27724),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__4800 (
            .O(N__27721),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__4799 (
            .O(N__27714),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__4798 (
            .O(N__27711),
            .I(N__27708));
    LocalMux I__4797 (
            .O(N__27708),
            .I(N__27704));
    InMux I__4796 (
            .O(N__27707),
            .I(N__27701));
    Span4Mux_v I__4795 (
            .O(N__27704),
            .I(N__27696));
    LocalMux I__4794 (
            .O(N__27701),
            .I(N__27696));
    Span4Mux_v I__4793 (
            .O(N__27696),
            .I(N__27692));
    InMux I__4792 (
            .O(N__27695),
            .I(N__27689));
    Odrv4 I__4791 (
            .O(N__27692),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__4790 (
            .O(N__27689),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__4789 (
            .O(N__27684),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__4788 (
            .O(N__27681),
            .I(N__27678));
    LocalMux I__4787 (
            .O(N__27678),
            .I(N__27675));
    Span4Mux_v I__4786 (
            .O(N__27675),
            .I(N__27672));
    Span4Mux_h I__4785 (
            .O(N__27672),
            .I(N__27669));
    Span4Mux_v I__4784 (
            .O(N__27669),
            .I(N__27666));
    Odrv4 I__4783 (
            .O(N__27666),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__4782 (
            .O(N__27663),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__4781 (
            .O(N__27660),
            .I(N__27657));
    LocalMux I__4780 (
            .O(N__27657),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__4779 (
            .O(N__27654),
            .I(N__27649));
    InMux I__4778 (
            .O(N__27653),
            .I(N__27646));
    InMux I__4777 (
            .O(N__27652),
            .I(N__27643));
    InMux I__4776 (
            .O(N__27649),
            .I(N__27640));
    LocalMux I__4775 (
            .O(N__27646),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__4774 (
            .O(N__27643),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__4773 (
            .O(N__27640),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__4772 (
            .O(N__27633),
            .I(N__27630));
    LocalMux I__4771 (
            .O(N__27630),
            .I(N__27627));
    Span4Mux_v I__4770 (
            .O(N__27627),
            .I(N__27622));
    InMux I__4769 (
            .O(N__27626),
            .I(N__27617));
    InMux I__4768 (
            .O(N__27625),
            .I(N__27617));
    Odrv4 I__4767 (
            .O(N__27622),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__4766 (
            .O(N__27617),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__4765 (
            .O(N__27612),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__4764 (
            .O(N__27609),
            .I(N__27606));
    LocalMux I__4763 (
            .O(N__27606),
            .I(N__27603));
    Span4Mux_v I__4762 (
            .O(N__27603),
            .I(N__27598));
    InMux I__4761 (
            .O(N__27602),
            .I(N__27593));
    InMux I__4760 (
            .O(N__27601),
            .I(N__27593));
    Odrv4 I__4759 (
            .O(N__27598),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__4758 (
            .O(N__27593),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__4757 (
            .O(N__27588),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__4756 (
            .O(N__27585),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    CascadeMux I__4755 (
            .O(N__27582),
            .I(N__27579));
    InMux I__4754 (
            .O(N__27579),
            .I(N__27576));
    LocalMux I__4753 (
            .O(N__27576),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__4752 (
            .O(N__27573),
            .I(N__27570));
    InMux I__4751 (
            .O(N__27570),
            .I(N__27567));
    LocalMux I__4750 (
            .O(N__27567),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__4749 (
            .O(N__27564),
            .I(N__27561));
    InMux I__4748 (
            .O(N__27561),
            .I(N__27558));
    LocalMux I__4747 (
            .O(N__27558),
            .I(N__27555));
    Odrv4 I__4746 (
            .O(N__27555),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__4745 (
            .O(N__27552),
            .I(N__27549));
    InMux I__4744 (
            .O(N__27549),
            .I(N__27546));
    LocalMux I__4743 (
            .O(N__27546),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__4742 (
            .O(N__27543),
            .I(N__27540));
    InMux I__4741 (
            .O(N__27540),
            .I(N__27537));
    LocalMux I__4740 (
            .O(N__27537),
            .I(N__27534));
    Odrv4 I__4739 (
            .O(N__27534),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__4738 (
            .O(N__27531),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__4737 (
            .O(N__27528),
            .I(N__27525));
    LocalMux I__4736 (
            .O(N__27525),
            .I(N__27522));
    Span4Mux_h I__4735 (
            .O(N__27522),
            .I(N__27519));
    Span4Mux_v I__4734 (
            .O(N__27519),
            .I(N__27516));
    Odrv4 I__4733 (
            .O(N__27516),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__4732 (
            .O(N__27513),
            .I(N__27510));
    InMux I__4731 (
            .O(N__27510),
            .I(N__27507));
    LocalMux I__4730 (
            .O(N__27507),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__4729 (
            .O(N__27504),
            .I(N__27501));
    LocalMux I__4728 (
            .O(N__27501),
            .I(N__27498));
    Span4Mux_h I__4727 (
            .O(N__27498),
            .I(N__27494));
    InMux I__4726 (
            .O(N__27497),
            .I(N__27491));
    Odrv4 I__4725 (
            .O(N__27494),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    LocalMux I__4724 (
            .O(N__27491),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__4723 (
            .O(N__27486),
            .I(N__27483));
    LocalMux I__4722 (
            .O(N__27483),
            .I(N__27480));
    Span4Mux_h I__4721 (
            .O(N__27480),
            .I(N__27477));
    Sp12to4 I__4720 (
            .O(N__27477),
            .I(N__27474));
    Span12Mux_s10_v I__4719 (
            .O(N__27474),
            .I(N__27469));
    CascadeMux I__4718 (
            .O(N__27473),
            .I(N__27466));
    CascadeMux I__4717 (
            .O(N__27472),
            .I(N__27463));
    Span12Mux_v I__4716 (
            .O(N__27469),
            .I(N__27459));
    InMux I__4715 (
            .O(N__27466),
            .I(N__27456));
    InMux I__4714 (
            .O(N__27463),
            .I(N__27453));
    InMux I__4713 (
            .O(N__27462),
            .I(N__27450));
    Odrv12 I__4712 (
            .O(N__27459),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__4711 (
            .O(N__27456),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__4710 (
            .O(N__27453),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__4709 (
            .O(N__27450),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__4708 (
            .O(N__27441),
            .I(N__27436));
    InMux I__4707 (
            .O(N__27440),
            .I(N__27433));
    InMux I__4706 (
            .O(N__27439),
            .I(N__27430));
    LocalMux I__4705 (
            .O(N__27436),
            .I(N__27427));
    LocalMux I__4704 (
            .O(N__27433),
            .I(N__27424));
    LocalMux I__4703 (
            .O(N__27430),
            .I(N__27421));
    Span4Mux_v I__4702 (
            .O(N__27427),
            .I(N__27418));
    Span4Mux_h I__4701 (
            .O(N__27424),
            .I(N__27415));
    Odrv4 I__4700 (
            .O(N__27421),
            .I(il_max_comp2_D2));
    Odrv4 I__4699 (
            .O(N__27418),
            .I(il_max_comp2_D2));
    Odrv4 I__4698 (
            .O(N__27415),
            .I(il_max_comp2_D2));
    CascadeMux I__4697 (
            .O(N__27408),
            .I(N__27405));
    InMux I__4696 (
            .O(N__27405),
            .I(N__27402));
    LocalMux I__4695 (
            .O(N__27402),
            .I(N__27399));
    Span4Mux_h I__4694 (
            .O(N__27399),
            .I(N__27396));
    Odrv4 I__4693 (
            .O(N__27396),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__4692 (
            .O(N__27393),
            .I(N__27390));
    InMux I__4691 (
            .O(N__27390),
            .I(N__27387));
    LocalMux I__4690 (
            .O(N__27387),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__4689 (
            .O(N__27384),
            .I(N__27381));
    InMux I__4688 (
            .O(N__27381),
            .I(N__27378));
    LocalMux I__4687 (
            .O(N__27378),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__4686 (
            .O(N__27375),
            .I(N__27372));
    InMux I__4685 (
            .O(N__27372),
            .I(N__27369));
    LocalMux I__4684 (
            .O(N__27369),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__4683 (
            .O(N__27366),
            .I(N__27363));
    InMux I__4682 (
            .O(N__27363),
            .I(N__27360));
    LocalMux I__4681 (
            .O(N__27360),
            .I(N__27357));
    Odrv4 I__4680 (
            .O(N__27357),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__4679 (
            .O(N__27354),
            .I(N__27351));
    LocalMux I__4678 (
            .O(N__27351),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__4677 (
            .O(N__27348),
            .I(N__27345));
    LocalMux I__4676 (
            .O(N__27345),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__4675 (
            .O(N__27342),
            .I(N__27339));
    LocalMux I__4674 (
            .O(N__27339),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__4673 (
            .O(N__27336),
            .I(N__27333));
    LocalMux I__4672 (
            .O(N__27333),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    InMux I__4671 (
            .O(N__27330),
            .I(N__27327));
    LocalMux I__4670 (
            .O(N__27327),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__4669 (
            .O(N__27324),
            .I(N__27321));
    LocalMux I__4668 (
            .O(N__27321),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__4667 (
            .O(N__27318),
            .I(N__27315));
    LocalMux I__4666 (
            .O(N__27315),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__4665 (
            .O(N__27312),
            .I(N__27309));
    LocalMux I__4664 (
            .O(N__27309),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__4663 (
            .O(N__27306),
            .I(N__27303));
    LocalMux I__4662 (
            .O(N__27303),
            .I(N__27300));
    Odrv4 I__4661 (
            .O(N__27300),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__4660 (
            .O(N__27297),
            .I(N__27294));
    LocalMux I__4659 (
            .O(N__27294),
            .I(N__27291));
    Span4Mux_h I__4658 (
            .O(N__27291),
            .I(N__27288));
    Odrv4 I__4657 (
            .O(N__27288),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__4656 (
            .O(N__27285),
            .I(N__27282));
    LocalMux I__4655 (
            .O(N__27282),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    InMux I__4654 (
            .O(N__27279),
            .I(N__27276));
    LocalMux I__4653 (
            .O(N__27276),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    InMux I__4652 (
            .O(N__27273),
            .I(N__27270));
    LocalMux I__4651 (
            .O(N__27270),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    InMux I__4650 (
            .O(N__27267),
            .I(N__27264));
    LocalMux I__4649 (
            .O(N__27264),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__4648 (
            .O(N__27261),
            .I(N__27258));
    LocalMux I__4647 (
            .O(N__27258),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__4646 (
            .O(N__27255),
            .I(N__27252));
    LocalMux I__4645 (
            .O(N__27252),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__4644 (
            .O(N__27249),
            .I(N__27246));
    LocalMux I__4643 (
            .O(N__27246),
            .I(N__27243));
    Odrv4 I__4642 (
            .O(N__27243),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__4641 (
            .O(N__27240),
            .I(N__27237));
    LocalMux I__4640 (
            .O(N__27237),
            .I(N__27234));
    Odrv4 I__4639 (
            .O(N__27234),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__4638 (
            .O(N__27231),
            .I(N__27228));
    LocalMux I__4637 (
            .O(N__27228),
            .I(N__27225));
    Span4Mux_v I__4636 (
            .O(N__27225),
            .I(N__27222));
    Odrv4 I__4635 (
            .O(N__27222),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__4634 (
            .O(N__27219),
            .I(N__27216));
    LocalMux I__4633 (
            .O(N__27216),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    CascadeMux I__4632 (
            .O(N__27213),
            .I(N__27210));
    InMux I__4631 (
            .O(N__27210),
            .I(N__27207));
    LocalMux I__4630 (
            .O(N__27207),
            .I(N__27204));
    Span4Mux_v I__4629 (
            .O(N__27204),
            .I(N__27201));
    Odrv4 I__4628 (
            .O(N__27201),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__4627 (
            .O(N__27198),
            .I(N__27195));
    LocalMux I__4626 (
            .O(N__27195),
            .I(N__27192));
    Span4Mux_v I__4625 (
            .O(N__27192),
            .I(N__27189));
    Odrv4 I__4624 (
            .O(N__27189),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__4623 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__4622 (
            .O(N__27183),
            .I(N__27180));
    Span4Mux_v I__4621 (
            .O(N__27180),
            .I(N__27177));
    Odrv4 I__4620 (
            .O(N__27177),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__4619 (
            .O(N__27174),
            .I(N__27171));
    LocalMux I__4618 (
            .O(N__27171),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__4617 (
            .O(N__27168),
            .I(N__27165));
    InMux I__4616 (
            .O(N__27165),
            .I(N__27162));
    LocalMux I__4615 (
            .O(N__27162),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    InMux I__4614 (
            .O(N__27159),
            .I(N__27156));
    LocalMux I__4613 (
            .O(N__27156),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__4612 (
            .O(N__27153),
            .I(N__27150));
    InMux I__4611 (
            .O(N__27150),
            .I(N__27147));
    LocalMux I__4610 (
            .O(N__27147),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    CascadeMux I__4609 (
            .O(N__27144),
            .I(N__27141));
    InMux I__4608 (
            .O(N__27141),
            .I(N__27138));
    LocalMux I__4607 (
            .O(N__27138),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__4606 (
            .O(N__27135),
            .I(N__27132));
    LocalMux I__4605 (
            .O(N__27132),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__4604 (
            .O(N__27129),
            .I(N__27126));
    LocalMux I__4603 (
            .O(N__27126),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__4602 (
            .O(N__27123),
            .I(N__27120));
    LocalMux I__4601 (
            .O(N__27120),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__4600 (
            .O(N__27117),
            .I(N__27114));
    LocalMux I__4599 (
            .O(N__27114),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__4598 (
            .O(N__27111),
            .I(N__27108));
    LocalMux I__4597 (
            .O(N__27108),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__4596 (
            .O(N__27105),
            .I(N__27102));
    LocalMux I__4595 (
            .O(N__27102),
            .I(N__27099));
    Span4Mux_v I__4594 (
            .O(N__27099),
            .I(N__27096));
    Odrv4 I__4593 (
            .O(N__27096),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__4592 (
            .O(N__27093),
            .I(N__27074));
    InMux I__4591 (
            .O(N__27092),
            .I(N__27071));
    InMux I__4590 (
            .O(N__27091),
            .I(N__27054));
    InMux I__4589 (
            .O(N__27090),
            .I(N__27054));
    InMux I__4588 (
            .O(N__27089),
            .I(N__27054));
    InMux I__4587 (
            .O(N__27088),
            .I(N__27054));
    InMux I__4586 (
            .O(N__27087),
            .I(N__27054));
    InMux I__4585 (
            .O(N__27086),
            .I(N__27054));
    InMux I__4584 (
            .O(N__27085),
            .I(N__27054));
    InMux I__4583 (
            .O(N__27084),
            .I(N__27054));
    InMux I__4582 (
            .O(N__27083),
            .I(N__27041));
    InMux I__4581 (
            .O(N__27082),
            .I(N__27041));
    InMux I__4580 (
            .O(N__27081),
            .I(N__27041));
    InMux I__4579 (
            .O(N__27080),
            .I(N__27041));
    InMux I__4578 (
            .O(N__27079),
            .I(N__27041));
    InMux I__4577 (
            .O(N__27078),
            .I(N__27041));
    InMux I__4576 (
            .O(N__27077),
            .I(N__27038));
    LocalMux I__4575 (
            .O(N__27074),
            .I(N__27033));
    LocalMux I__4574 (
            .O(N__27071),
            .I(N__27033));
    LocalMux I__4573 (
            .O(N__27054),
            .I(N__27030));
    LocalMux I__4572 (
            .O(N__27041),
            .I(N__27027));
    LocalMux I__4571 (
            .O(N__27038),
            .I(N__27014));
    Span4Mux_v I__4570 (
            .O(N__27033),
            .I(N__27011));
    Span4Mux_v I__4569 (
            .O(N__27030),
            .I(N__27006));
    Span4Mux_v I__4568 (
            .O(N__27027),
            .I(N__27006));
    InMux I__4567 (
            .O(N__27026),
            .I(N__26997));
    InMux I__4566 (
            .O(N__27025),
            .I(N__26997));
    InMux I__4565 (
            .O(N__27024),
            .I(N__26997));
    InMux I__4564 (
            .O(N__27023),
            .I(N__26997));
    InMux I__4563 (
            .O(N__27022),
            .I(N__26986));
    InMux I__4562 (
            .O(N__27021),
            .I(N__26986));
    InMux I__4561 (
            .O(N__27020),
            .I(N__26986));
    InMux I__4560 (
            .O(N__27019),
            .I(N__26986));
    InMux I__4559 (
            .O(N__27018),
            .I(N__26986));
    InMux I__4558 (
            .O(N__27017),
            .I(N__26983));
    Odrv4 I__4557 (
            .O(N__27014),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__4556 (
            .O(N__27011),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__4555 (
            .O(N__27006),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__4554 (
            .O(N__26997),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__4553 (
            .O(N__26986),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__4552 (
            .O(N__26983),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    CascadeMux I__4551 (
            .O(N__26970),
            .I(N__26966));
    InMux I__4550 (
            .O(N__26969),
            .I(N__26963));
    InMux I__4549 (
            .O(N__26966),
            .I(N__26960));
    LocalMux I__4548 (
            .O(N__26963),
            .I(N__26955));
    LocalMux I__4547 (
            .O(N__26960),
            .I(N__26955));
    Span12Mux_v I__4546 (
            .O(N__26955),
            .I(N__26952));
    Odrv12 I__4545 (
            .O(N__26952),
            .I(\current_shift_inst.N_1819_i ));
    InMux I__4544 (
            .O(N__26949),
            .I(N__26946));
    LocalMux I__4543 (
            .O(N__26946),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__4542 (
            .O(N__26943),
            .I(N__26940));
    InMux I__4541 (
            .O(N__26940),
            .I(N__26937));
    LocalMux I__4540 (
            .O(N__26937),
            .I(N__26934));
    Span4Mux_v I__4539 (
            .O(N__26934),
            .I(N__26931));
    Odrv4 I__4538 (
            .O(N__26931),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    InMux I__4537 (
            .O(N__26928),
            .I(N__26925));
    LocalMux I__4536 (
            .O(N__26925),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    InMux I__4535 (
            .O(N__26922),
            .I(N__26919));
    LocalMux I__4534 (
            .O(N__26919),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__4533 (
            .O(N__26916),
            .I(N__26913));
    LocalMux I__4532 (
            .O(N__26913),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__4531 (
            .O(N__26910),
            .I(N__26907));
    LocalMux I__4530 (
            .O(N__26907),
            .I(N__26904));
    Span4Mux_v I__4529 (
            .O(N__26904),
            .I(N__26901));
    Odrv4 I__4528 (
            .O(N__26901),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    InMux I__4527 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__4526 (
            .O(N__26895),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__4525 (
            .O(N__26892),
            .I(N__26889));
    LocalMux I__4524 (
            .O(N__26889),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__4523 (
            .O(N__26886),
            .I(N__26883));
    InMux I__4522 (
            .O(N__26883),
            .I(N__26880));
    LocalMux I__4521 (
            .O(N__26880),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__4520 (
            .O(N__26877),
            .I(N__26874));
    LocalMux I__4519 (
            .O(N__26874),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__4518 (
            .O(N__26871),
            .I(N__26868));
    LocalMux I__4517 (
            .O(N__26868),
            .I(N__26865));
    Span12Mux_v I__4516 (
            .O(N__26865),
            .I(N__26862));
    Odrv12 I__4515 (
            .O(N__26862),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__4514 (
            .O(N__26859),
            .I(N__26856));
    LocalMux I__4513 (
            .O(N__26856),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__4512 (
            .O(N__26853),
            .I(N__26850));
    LocalMux I__4511 (
            .O(N__26850),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__4510 (
            .O(N__26847),
            .I(N__26844));
    LocalMux I__4509 (
            .O(N__26844),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__4508 (
            .O(N__26841),
            .I(N__26838));
    LocalMux I__4507 (
            .O(N__26838),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__4506 (
            .O(N__26835),
            .I(N__26832));
    LocalMux I__4505 (
            .O(N__26832),
            .I(N__26829));
    Span4Mux_v I__4504 (
            .O(N__26829),
            .I(N__26826));
    Odrv4 I__4503 (
            .O(N__26826),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__4502 (
            .O(N__26823),
            .I(N__26820));
    LocalMux I__4501 (
            .O(N__26820),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__4500 (
            .O(N__26817),
            .I(N__26814));
    LocalMux I__4499 (
            .O(N__26814),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__4498 (
            .O(N__26811),
            .I(N__26808));
    LocalMux I__4497 (
            .O(N__26808),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__4496 (
            .O(N__26805),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__4495 (
            .O(N__26802),
            .I(N__26799));
    InMux I__4494 (
            .O(N__26799),
            .I(N__26796));
    LocalMux I__4493 (
            .O(N__26796),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__4492 (
            .O(N__26793),
            .I(N__26790));
    InMux I__4491 (
            .O(N__26790),
            .I(N__26787));
    LocalMux I__4490 (
            .O(N__26787),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__4489 (
            .O(N__26784),
            .I(N__26781));
    InMux I__4488 (
            .O(N__26781),
            .I(N__26778));
    LocalMux I__4487 (
            .O(N__26778),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__4486 (
            .O(N__26775),
            .I(N__26772));
    LocalMux I__4485 (
            .O(N__26772),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__4484 (
            .O(N__26769),
            .I(N__26766));
    InMux I__4483 (
            .O(N__26766),
            .I(N__26763));
    LocalMux I__4482 (
            .O(N__26763),
            .I(N__26759));
    CascadeMux I__4481 (
            .O(N__26762),
            .I(N__26756));
    Span4Mux_v I__4480 (
            .O(N__26759),
            .I(N__26751));
    InMux I__4479 (
            .O(N__26756),
            .I(N__26748));
    CascadeMux I__4478 (
            .O(N__26755),
            .I(N__26745));
    CascadeMux I__4477 (
            .O(N__26754),
            .I(N__26742));
    Span4Mux_v I__4476 (
            .O(N__26751),
            .I(N__26739));
    LocalMux I__4475 (
            .O(N__26748),
            .I(N__26736));
    InMux I__4474 (
            .O(N__26745),
            .I(N__26733));
    InMux I__4473 (
            .O(N__26742),
            .I(N__26730));
    Odrv4 I__4472 (
            .O(N__26739),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__4471 (
            .O(N__26736),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__4470 (
            .O(N__26733),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__4469 (
            .O(N__26730),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__4468 (
            .O(N__26721),
            .I(N__26718));
    LocalMux I__4467 (
            .O(N__26718),
            .I(N__26715));
    Span4Mux_v I__4466 (
            .O(N__26715),
            .I(N__26712));
    Odrv4 I__4465 (
            .O(N__26712),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__4464 (
            .O(N__26709),
            .I(N__26706));
    LocalMux I__4463 (
            .O(N__26706),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__4462 (
            .O(N__26703),
            .I(N__26700));
    LocalMux I__4461 (
            .O(N__26700),
            .I(N__26697));
    Span4Mux_v I__4460 (
            .O(N__26697),
            .I(N__26691));
    InMux I__4459 (
            .O(N__26696),
            .I(N__26684));
    InMux I__4458 (
            .O(N__26695),
            .I(N__26684));
    InMux I__4457 (
            .O(N__26694),
            .I(N__26684));
    Odrv4 I__4456 (
            .O(N__26691),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__4455 (
            .O(N__26684),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__4454 (
            .O(N__26679),
            .I(N__26676));
    LocalMux I__4453 (
            .O(N__26676),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__4452 (
            .O(N__26673),
            .I(N__26670));
    LocalMux I__4451 (
            .O(N__26670),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__4450 (
            .O(N__26667),
            .I(N__26664));
    InMux I__4449 (
            .O(N__26664),
            .I(N__26661));
    LocalMux I__4448 (
            .O(N__26661),
            .I(N__26658));
    Odrv4 I__4447 (
            .O(N__26658),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__4446 (
            .O(N__26655),
            .I(N__26651));
    InMux I__4445 (
            .O(N__26654),
            .I(N__26648));
    LocalMux I__4444 (
            .O(N__26651),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__4443 (
            .O(N__26648),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__4442 (
            .O(N__26643),
            .I(N__26640));
    LocalMux I__4441 (
            .O(N__26640),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__4440 (
            .O(N__26637),
            .I(N__26633));
    InMux I__4439 (
            .O(N__26636),
            .I(N__26630));
    LocalMux I__4438 (
            .O(N__26633),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__4437 (
            .O(N__26630),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__4436 (
            .O(N__26625),
            .I(N__26622));
    LocalMux I__4435 (
            .O(N__26622),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__4434 (
            .O(N__26619),
            .I(N__26615));
    InMux I__4433 (
            .O(N__26618),
            .I(N__26612));
    LocalMux I__4432 (
            .O(N__26615),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__4431 (
            .O(N__26612),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__4430 (
            .O(N__26607),
            .I(N__26604));
    LocalMux I__4429 (
            .O(N__26604),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__4428 (
            .O(N__26601),
            .I(N__26598));
    InMux I__4427 (
            .O(N__26598),
            .I(N__26595));
    LocalMux I__4426 (
            .O(N__26595),
            .I(N__26592));
    Odrv12 I__4425 (
            .O(N__26592),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    InMux I__4424 (
            .O(N__26589),
            .I(N__26586));
    LocalMux I__4423 (
            .O(N__26586),
            .I(N__26582));
    InMux I__4422 (
            .O(N__26585),
            .I(N__26579));
    Span4Mux_h I__4421 (
            .O(N__26582),
            .I(N__26576));
    LocalMux I__4420 (
            .O(N__26579),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__4419 (
            .O(N__26576),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__4418 (
            .O(N__26571),
            .I(N__26568));
    LocalMux I__4417 (
            .O(N__26568),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ));
    InMux I__4416 (
            .O(N__26565),
            .I(N__26561));
    InMux I__4415 (
            .O(N__26564),
            .I(N__26558));
    LocalMux I__4414 (
            .O(N__26561),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__4413 (
            .O(N__26558),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__4412 (
            .O(N__26553),
            .I(N__26550));
    LocalMux I__4411 (
            .O(N__26550),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ));
    InMux I__4410 (
            .O(N__26547),
            .I(N__26543));
    InMux I__4409 (
            .O(N__26546),
            .I(N__26540));
    LocalMux I__4408 (
            .O(N__26543),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__4407 (
            .O(N__26540),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__4406 (
            .O(N__26535),
            .I(N__26532));
    LocalMux I__4405 (
            .O(N__26532),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ));
    InMux I__4404 (
            .O(N__26529),
            .I(N__26525));
    InMux I__4403 (
            .O(N__26528),
            .I(N__26522));
    LocalMux I__4402 (
            .O(N__26525),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__4401 (
            .O(N__26522),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__4400 (
            .O(N__26517),
            .I(N__26514));
    LocalMux I__4399 (
            .O(N__26514),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ));
    CascadeMux I__4398 (
            .O(N__26511),
            .I(N__26508));
    InMux I__4397 (
            .O(N__26508),
            .I(N__26505));
    LocalMux I__4396 (
            .O(N__26505),
            .I(N__26502));
    Odrv4 I__4395 (
            .O(N__26502),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__4394 (
            .O(N__26499),
            .I(N__26496));
    InMux I__4393 (
            .O(N__26496),
            .I(N__26492));
    InMux I__4392 (
            .O(N__26495),
            .I(N__26489));
    LocalMux I__4391 (
            .O(N__26492),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__4390 (
            .O(N__26489),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__4389 (
            .O(N__26484),
            .I(N__26481));
    LocalMux I__4388 (
            .O(N__26481),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__4387 (
            .O(N__26478),
            .I(N__26474));
    InMux I__4386 (
            .O(N__26477),
            .I(N__26471));
    LocalMux I__4385 (
            .O(N__26474),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__4384 (
            .O(N__26471),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__4383 (
            .O(N__26466),
            .I(N__26463));
    LocalMux I__4382 (
            .O(N__26463),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__4381 (
            .O(N__26460),
            .I(N__26456));
    InMux I__4380 (
            .O(N__26459),
            .I(N__26453));
    LocalMux I__4379 (
            .O(N__26456),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__4378 (
            .O(N__26453),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__4377 (
            .O(N__26448),
            .I(N__26445));
    InMux I__4376 (
            .O(N__26445),
            .I(N__26442));
    LocalMux I__4375 (
            .O(N__26442),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__4374 (
            .O(N__26439),
            .I(N__26436));
    LocalMux I__4373 (
            .O(N__26436),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__4372 (
            .O(N__26433),
            .I(N__26429));
    InMux I__4371 (
            .O(N__26432),
            .I(N__26426));
    LocalMux I__4370 (
            .O(N__26429),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__4369 (
            .O(N__26426),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__4368 (
            .O(N__26421),
            .I(N__26418));
    InMux I__4367 (
            .O(N__26418),
            .I(N__26415));
    LocalMux I__4366 (
            .O(N__26415),
            .I(N__26412));
    Odrv4 I__4365 (
            .O(N__26412),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    InMux I__4364 (
            .O(N__26409),
            .I(N__26406));
    LocalMux I__4363 (
            .O(N__26406),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__4362 (
            .O(N__26403),
            .I(N__26399));
    InMux I__4361 (
            .O(N__26402),
            .I(N__26396));
    LocalMux I__4360 (
            .O(N__26399),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__4359 (
            .O(N__26396),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__4358 (
            .O(N__26391),
            .I(N__26388));
    LocalMux I__4357 (
            .O(N__26388),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__4356 (
            .O(N__26385),
            .I(N__26381));
    InMux I__4355 (
            .O(N__26384),
            .I(N__26378));
    LocalMux I__4354 (
            .O(N__26381),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__4353 (
            .O(N__26378),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__4352 (
            .O(N__26373),
            .I(N__26370));
    LocalMux I__4351 (
            .O(N__26370),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__4350 (
            .O(N__26367),
            .I(N__26364));
    InMux I__4349 (
            .O(N__26364),
            .I(N__26361));
    LocalMux I__4348 (
            .O(N__26361),
            .I(N__26358));
    Span4Mux_h I__4347 (
            .O(N__26358),
            .I(N__26355));
    Odrv4 I__4346 (
            .O(N__26355),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__4345 (
            .O(N__26352),
            .I(N__26348));
    InMux I__4344 (
            .O(N__26351),
            .I(N__26345));
    LocalMux I__4343 (
            .O(N__26348),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__4342 (
            .O(N__26345),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__4341 (
            .O(N__26340),
            .I(N__26337));
    LocalMux I__4340 (
            .O(N__26337),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__4339 (
            .O(N__26334),
            .I(N__26330));
    InMux I__4338 (
            .O(N__26333),
            .I(N__26327));
    LocalMux I__4337 (
            .O(N__26330),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__4336 (
            .O(N__26327),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__4335 (
            .O(N__26322),
            .I(N__26319));
    LocalMux I__4334 (
            .O(N__26319),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__4333 (
            .O(N__26316),
            .I(N__26312));
    InMux I__4332 (
            .O(N__26315),
            .I(N__26308));
    InMux I__4331 (
            .O(N__26312),
            .I(N__26305));
    InMux I__4330 (
            .O(N__26311),
            .I(N__26302));
    LocalMux I__4329 (
            .O(N__26308),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__4328 (
            .O(N__26305),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__4327 (
            .O(N__26302),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__4326 (
            .O(N__26295),
            .I(N__26292));
    LocalMux I__4325 (
            .O(N__26292),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__4324 (
            .O(N__26289),
            .I(N__26285));
    InMux I__4323 (
            .O(N__26288),
            .I(N__26282));
    LocalMux I__4322 (
            .O(N__26285),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__4321 (
            .O(N__26282),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__4320 (
            .O(N__26277),
            .I(N__26274));
    LocalMux I__4319 (
            .O(N__26274),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__4318 (
            .O(N__26271),
            .I(N__26268));
    InMux I__4317 (
            .O(N__26268),
            .I(N__26264));
    InMux I__4316 (
            .O(N__26267),
            .I(N__26261));
    LocalMux I__4315 (
            .O(N__26264),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__4314 (
            .O(N__26261),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__4313 (
            .O(N__26256),
            .I(N__26253));
    LocalMux I__4312 (
            .O(N__26253),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__4311 (
            .O(N__26250),
            .I(N__26246));
    InMux I__4310 (
            .O(N__26249),
            .I(N__26243));
    LocalMux I__4309 (
            .O(N__26246),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__4308 (
            .O(N__26243),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__4307 (
            .O(N__26238),
            .I(N__26235));
    LocalMux I__4306 (
            .O(N__26235),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__4305 (
            .O(N__26232),
            .I(N__26229));
    LocalMux I__4304 (
            .O(N__26229),
            .I(N__26226));
    Span4Mux_v I__4303 (
            .O(N__26226),
            .I(N__26223));
    Odrv4 I__4302 (
            .O(N__26223),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__4301 (
            .O(N__26220),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__4300 (
            .O(N__26217),
            .I(N__26214));
    LocalMux I__4299 (
            .O(N__26214),
            .I(N__26211));
    Sp12to4 I__4298 (
            .O(N__26211),
            .I(N__26208));
    Odrv12 I__4297 (
            .O(N__26208),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__4296 (
            .O(N__26205),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__4295 (
            .O(N__26202),
            .I(N__26199));
    LocalMux I__4294 (
            .O(N__26199),
            .I(N__26196));
    Sp12to4 I__4293 (
            .O(N__26196),
            .I(N__26193));
    Odrv12 I__4292 (
            .O(N__26193),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__4291 (
            .O(N__26190),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__4290 (
            .O(N__26187),
            .I(N__26184));
    LocalMux I__4289 (
            .O(N__26184),
            .I(N__26181));
    Odrv4 I__4288 (
            .O(N__26181),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__4287 (
            .O(N__26178),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__4286 (
            .O(N__26175),
            .I(N__26172));
    LocalMux I__4285 (
            .O(N__26172),
            .I(N__26169));
    Span4Mux_v I__4284 (
            .O(N__26169),
            .I(N__26166));
    Odrv4 I__4283 (
            .O(N__26166),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__4282 (
            .O(N__26163),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__4281 (
            .O(N__26160),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    CascadeMux I__4280 (
            .O(N__26157),
            .I(N__26154));
    InMux I__4279 (
            .O(N__26154),
            .I(N__26151));
    LocalMux I__4278 (
            .O(N__26151),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    IoInMux I__4277 (
            .O(N__26148),
            .I(N__26145));
    LocalMux I__4276 (
            .O(N__26145),
            .I(N__26142));
    Odrv12 I__4275 (
            .O(N__26142),
            .I(s3_phy_c));
    InMux I__4274 (
            .O(N__26139),
            .I(N__26136));
    LocalMux I__4273 (
            .O(N__26136),
            .I(N__26133));
    Span4Mux_v I__4272 (
            .O(N__26133),
            .I(N__26130));
    Odrv4 I__4271 (
            .O(N__26130),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__4270 (
            .O(N__26127),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__4269 (
            .O(N__26124),
            .I(N__26121));
    LocalMux I__4268 (
            .O(N__26121),
            .I(N__26118));
    Span4Mux_v I__4267 (
            .O(N__26118),
            .I(N__26115));
    Odrv4 I__4266 (
            .O(N__26115),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__4265 (
            .O(N__26112),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__4264 (
            .O(N__26109),
            .I(N__26106));
    LocalMux I__4263 (
            .O(N__26106),
            .I(N__26103));
    Span4Mux_v I__4262 (
            .O(N__26103),
            .I(N__26100));
    Span4Mux_h I__4261 (
            .O(N__26100),
            .I(N__26097));
    Odrv4 I__4260 (
            .O(N__26097),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__4259 (
            .O(N__26094),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    InMux I__4258 (
            .O(N__26091),
            .I(N__26088));
    LocalMux I__4257 (
            .O(N__26088),
            .I(N__26085));
    Span4Mux_v I__4256 (
            .O(N__26085),
            .I(N__26082));
    Odrv4 I__4255 (
            .O(N__26082),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__4254 (
            .O(N__26079),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__4253 (
            .O(N__26076),
            .I(N__26073));
    LocalMux I__4252 (
            .O(N__26073),
            .I(N__26070));
    Span4Mux_v I__4251 (
            .O(N__26070),
            .I(N__26067));
    Odrv4 I__4250 (
            .O(N__26067),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__4249 (
            .O(N__26064),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__4248 (
            .O(N__26061),
            .I(N__26058));
    LocalMux I__4247 (
            .O(N__26058),
            .I(N__26055));
    Span4Mux_v I__4246 (
            .O(N__26055),
            .I(N__26052));
    Odrv4 I__4245 (
            .O(N__26052),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__4244 (
            .O(N__26049),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__4243 (
            .O(N__26046),
            .I(N__26043));
    LocalMux I__4242 (
            .O(N__26043),
            .I(N__26040));
    Span4Mux_h I__4241 (
            .O(N__26040),
            .I(N__26037));
    Odrv4 I__4240 (
            .O(N__26037),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__4239 (
            .O(N__26034),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__4238 (
            .O(N__26031),
            .I(N__26028));
    LocalMux I__4237 (
            .O(N__26028),
            .I(N__26025));
    Span4Mux_v I__4236 (
            .O(N__26025),
            .I(N__26022));
    Odrv4 I__4235 (
            .O(N__26022),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__4234 (
            .O(N__26019),
            .I(bfn_9_22_0_));
    InMux I__4233 (
            .O(N__26016),
            .I(N__26013));
    LocalMux I__4232 (
            .O(N__26013),
            .I(N__26010));
    Span4Mux_v I__4231 (
            .O(N__26010),
            .I(N__26007));
    Odrv4 I__4230 (
            .O(N__26007),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__4229 (
            .O(N__26004),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__4228 (
            .O(N__26001),
            .I(N__25998));
    LocalMux I__4227 (
            .O(N__25998),
            .I(N__25995));
    Odrv12 I__4226 (
            .O(N__25995),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__4225 (
            .O(N__25992),
            .I(N__25989));
    LocalMux I__4224 (
            .O(N__25989),
            .I(N__25986));
    Span4Mux_v I__4223 (
            .O(N__25986),
            .I(N__25983));
    Odrv4 I__4222 (
            .O(N__25983),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__4221 (
            .O(N__25980),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__4220 (
            .O(N__25977),
            .I(N__25974));
    LocalMux I__4219 (
            .O(N__25974),
            .I(N__25971));
    Odrv4 I__4218 (
            .O(N__25971),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__4217 (
            .O(N__25968),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__4216 (
            .O(N__25965),
            .I(N__25962));
    LocalMux I__4215 (
            .O(N__25962),
            .I(N__25959));
    Span4Mux_v I__4214 (
            .O(N__25959),
            .I(N__25956));
    Odrv4 I__4213 (
            .O(N__25956),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__4212 (
            .O(N__25953),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__4211 (
            .O(N__25950),
            .I(N__25947));
    LocalMux I__4210 (
            .O(N__25947),
            .I(N__25944));
    Span4Mux_v I__4209 (
            .O(N__25944),
            .I(N__25941));
    Odrv4 I__4208 (
            .O(N__25941),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__4207 (
            .O(N__25938),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__4206 (
            .O(N__25935),
            .I(N__25932));
    LocalMux I__4205 (
            .O(N__25932),
            .I(N__25929));
    Odrv4 I__4204 (
            .O(N__25929),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__4203 (
            .O(N__25926),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__4202 (
            .O(N__25923),
            .I(N__25920));
    LocalMux I__4201 (
            .O(N__25920),
            .I(N__25917));
    Span4Mux_h I__4200 (
            .O(N__25917),
            .I(N__25914));
    Span4Mux_v I__4199 (
            .O(N__25914),
            .I(N__25911));
    Odrv4 I__4198 (
            .O(N__25911),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__4197 (
            .O(N__25908),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__4196 (
            .O(N__25905),
            .I(N__25902));
    LocalMux I__4195 (
            .O(N__25902),
            .I(N__25899));
    Span4Mux_h I__4194 (
            .O(N__25899),
            .I(N__25896));
    Odrv4 I__4193 (
            .O(N__25896),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__4192 (
            .O(N__25893),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__4191 (
            .O(N__25890),
            .I(N__25887));
    LocalMux I__4190 (
            .O(N__25887),
            .I(N__25884));
    Span4Mux_v I__4189 (
            .O(N__25884),
            .I(N__25881));
    Odrv4 I__4188 (
            .O(N__25881),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__4187 (
            .O(N__25878),
            .I(bfn_9_21_0_));
    InMux I__4186 (
            .O(N__25875),
            .I(N__25872));
    LocalMux I__4185 (
            .O(N__25872),
            .I(N__25869));
    Span4Mux_h I__4184 (
            .O(N__25869),
            .I(N__25866));
    Odrv4 I__4183 (
            .O(N__25866),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__4182 (
            .O(N__25863),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__4181 (
            .O(N__25860),
            .I(N__25857));
    LocalMux I__4180 (
            .O(N__25857),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__4179 (
            .O(N__25854),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__4178 (
            .O(N__25851),
            .I(N__25848));
    LocalMux I__4177 (
            .O(N__25848),
            .I(N__25845));
    Span4Mux_v I__4176 (
            .O(N__25845),
            .I(N__25842));
    Odrv4 I__4175 (
            .O(N__25842),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__4174 (
            .O(N__25839),
            .I(bfn_9_20_0_));
    InMux I__4173 (
            .O(N__25836),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__4172 (
            .O(N__25833),
            .I(N__25830));
    LocalMux I__4171 (
            .O(N__25830),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ));
    InMux I__4170 (
            .O(N__25827),
            .I(N__25824));
    LocalMux I__4169 (
            .O(N__25824),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ));
    CascadeMux I__4168 (
            .O(N__25821),
            .I(N__25818));
    InMux I__4167 (
            .O(N__25818),
            .I(N__25815));
    LocalMux I__4166 (
            .O(N__25815),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ));
    InMux I__4165 (
            .O(N__25812),
            .I(N__25809));
    LocalMux I__4164 (
            .O(N__25809),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ));
    CascadeMux I__4163 (
            .O(N__25806),
            .I(N__25803));
    InMux I__4162 (
            .O(N__25803),
            .I(N__25800));
    LocalMux I__4161 (
            .O(N__25800),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ));
    InMux I__4160 (
            .O(N__25797),
            .I(N__25794));
    LocalMux I__4159 (
            .O(N__25794),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ));
    InMux I__4158 (
            .O(N__25791),
            .I(N__25788));
    LocalMux I__4157 (
            .O(N__25788),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ));
    InMux I__4156 (
            .O(N__25785),
            .I(N__25782));
    LocalMux I__4155 (
            .O(N__25782),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ));
    InMux I__4154 (
            .O(N__25779),
            .I(N__25776));
    LocalMux I__4153 (
            .O(N__25776),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ));
    InMux I__4152 (
            .O(N__25773),
            .I(N__25770));
    LocalMux I__4151 (
            .O(N__25770),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ));
    InMux I__4150 (
            .O(N__25767),
            .I(N__25764));
    LocalMux I__4149 (
            .O(N__25764),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ));
    InMux I__4148 (
            .O(N__25761),
            .I(N__25758));
    LocalMux I__4147 (
            .O(N__25758),
            .I(N__25755));
    Span4Mux_h I__4146 (
            .O(N__25755),
            .I(N__25752));
    Odrv4 I__4145 (
            .O(N__25752),
            .I(il_max_comp2_D1));
    InMux I__4144 (
            .O(N__25749),
            .I(N__25746));
    LocalMux I__4143 (
            .O(N__25746),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ));
    CascadeMux I__4142 (
            .O(N__25743),
            .I(N__25740));
    InMux I__4141 (
            .O(N__25740),
            .I(N__25737));
    LocalMux I__4140 (
            .O(N__25737),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ));
    InMux I__4139 (
            .O(N__25734),
            .I(N__25731));
    LocalMux I__4138 (
            .O(N__25731),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ));
    InMux I__4137 (
            .O(N__25728),
            .I(N__25725));
    LocalMux I__4136 (
            .O(N__25725),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ));
    CascadeMux I__4135 (
            .O(N__25722),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ));
    InMux I__4134 (
            .O(N__25719),
            .I(N__25716));
    LocalMux I__4133 (
            .O(N__25716),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ));
    InMux I__4132 (
            .O(N__25713),
            .I(N__25710));
    LocalMux I__4131 (
            .O(N__25710),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ));
    InMux I__4130 (
            .O(N__25707),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__4129 (
            .O(N__25704),
            .I(N__25701));
    LocalMux I__4128 (
            .O(N__25701),
            .I(N__25698));
    Span4Mux_v I__4127 (
            .O(N__25698),
            .I(N__25695));
    Odrv4 I__4126 (
            .O(N__25695),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__4125 (
            .O(N__25692),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__4124 (
            .O(N__25689),
            .I(N__25686));
    LocalMux I__4123 (
            .O(N__25686),
            .I(N__25683));
    Odrv12 I__4122 (
            .O(N__25683),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__4121 (
            .O(N__25680),
            .I(N__25677));
    LocalMux I__4120 (
            .O(N__25677),
            .I(N__25674));
    Odrv12 I__4119 (
            .O(N__25674),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__4118 (
            .O(N__25671),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__4117 (
            .O(N__25668),
            .I(N__25665));
    LocalMux I__4116 (
            .O(N__25665),
            .I(N__25662));
    Span4Mux_h I__4115 (
            .O(N__25662),
            .I(N__25659));
    Span4Mux_v I__4114 (
            .O(N__25659),
            .I(N__25656));
    Odrv4 I__4113 (
            .O(N__25656),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__4112 (
            .O(N__25653),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__4111 (
            .O(N__25650),
            .I(N__25647));
    LocalMux I__4110 (
            .O(N__25647),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__4109 (
            .O(N__25644),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__4108 (
            .O(N__25641),
            .I(N__25638));
    LocalMux I__4107 (
            .O(N__25638),
            .I(N__25635));
    Odrv12 I__4106 (
            .O(N__25635),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__4105 (
            .O(N__25632),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__4104 (
            .O(N__25629),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__4103 (
            .O(N__25626),
            .I(N__25623));
    LocalMux I__4102 (
            .O(N__25623),
            .I(N__25620));
    Span4Mux_h I__4101 (
            .O(N__25620),
            .I(N__25617));
    Span4Mux_v I__4100 (
            .O(N__25617),
            .I(N__25614));
    Odrv4 I__4099 (
            .O(N__25614),
            .I(\current_shift_inst.control_input_1_axb_25 ));
    IoInMux I__4098 (
            .O(N__25611),
            .I(N__25608));
    LocalMux I__4097 (
            .O(N__25608),
            .I(N__25605));
    Odrv12 I__4096 (
            .O(N__25605),
            .I(s4_phy_c));
    InMux I__4095 (
            .O(N__25602),
            .I(N__25599));
    LocalMux I__4094 (
            .O(N__25599),
            .I(N__25596));
    Odrv4 I__4093 (
            .O(N__25596),
            .I(il_max_comp1_D1));
    InMux I__4092 (
            .O(N__25593),
            .I(N__25590));
    LocalMux I__4091 (
            .O(N__25590),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__4090 (
            .O(N__25587),
            .I(N__25584));
    LocalMux I__4089 (
            .O(N__25584),
            .I(N__25581));
    Odrv12 I__4088 (
            .O(N__25581),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__4087 (
            .O(N__25578),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__4086 (
            .O(N__25575),
            .I(N__25572));
    LocalMux I__4085 (
            .O(N__25572),
            .I(N__25569));
    Odrv12 I__4084 (
            .O(N__25569),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__4083 (
            .O(N__25566),
            .I(N__25563));
    LocalMux I__4082 (
            .O(N__25563),
            .I(N__25560));
    Span4Mux_v I__4081 (
            .O(N__25560),
            .I(N__25557));
    Odrv4 I__4080 (
            .O(N__25557),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__4079 (
            .O(N__25554),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__4078 (
            .O(N__25551),
            .I(N__25548));
    LocalMux I__4077 (
            .O(N__25548),
            .I(N__25545));
    Odrv12 I__4076 (
            .O(N__25545),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__4075 (
            .O(N__25542),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    InMux I__4074 (
            .O(N__25539),
            .I(N__25536));
    LocalMux I__4073 (
            .O(N__25536),
            .I(N__25533));
    Odrv12 I__4072 (
            .O(N__25533),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__4071 (
            .O(N__25530),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__4070 (
            .O(N__25527),
            .I(N__25524));
    LocalMux I__4069 (
            .O(N__25524),
            .I(N__25521));
    Span4Mux_v I__4068 (
            .O(N__25521),
            .I(N__25518));
    Odrv4 I__4067 (
            .O(N__25518),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__4066 (
            .O(N__25515),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__4065 (
            .O(N__25512),
            .I(N__25509));
    LocalMux I__4064 (
            .O(N__25509),
            .I(N__25506));
    Span4Mux_h I__4063 (
            .O(N__25506),
            .I(N__25503));
    Span4Mux_v I__4062 (
            .O(N__25503),
            .I(N__25500));
    Odrv4 I__4061 (
            .O(N__25500),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__4060 (
            .O(N__25497),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__4059 (
            .O(N__25494),
            .I(N__25491));
    LocalMux I__4058 (
            .O(N__25491),
            .I(N__25488));
    Odrv12 I__4057 (
            .O(N__25488),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__4056 (
            .O(N__25485),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__4055 (
            .O(N__25482),
            .I(N__25479));
    LocalMux I__4054 (
            .O(N__25479),
            .I(N__25476));
    Span4Mux_v I__4053 (
            .O(N__25476),
            .I(N__25473));
    Odrv4 I__4052 (
            .O(N__25473),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__4051 (
            .O(N__25470),
            .I(bfn_8_22_0_));
    InMux I__4050 (
            .O(N__25467),
            .I(N__25464));
    LocalMux I__4049 (
            .O(N__25464),
            .I(N__25461));
    Span4Mux_v I__4048 (
            .O(N__25461),
            .I(N__25458));
    Odrv4 I__4047 (
            .O(N__25458),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__4046 (
            .O(N__25455),
            .I(N__25452));
    LocalMux I__4045 (
            .O(N__25452),
            .I(N__25449));
    Odrv12 I__4044 (
            .O(N__25449),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__4043 (
            .O(N__25446),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__4042 (
            .O(N__25443),
            .I(N__25440));
    LocalMux I__4041 (
            .O(N__25440),
            .I(N__25437));
    Odrv4 I__4040 (
            .O(N__25437),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__4039 (
            .O(N__25434),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__4038 (
            .O(N__25431),
            .I(N__25428));
    LocalMux I__4037 (
            .O(N__25428),
            .I(N__25425));
    Odrv12 I__4036 (
            .O(N__25425),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__4035 (
            .O(N__25422),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__4034 (
            .O(N__25419),
            .I(N__25416));
    LocalMux I__4033 (
            .O(N__25416),
            .I(N__25413));
    Odrv12 I__4032 (
            .O(N__25413),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__4031 (
            .O(N__25410),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__4030 (
            .O(N__25407),
            .I(N__25404));
    LocalMux I__4029 (
            .O(N__25404),
            .I(N__25401));
    Odrv4 I__4028 (
            .O(N__25401),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__4027 (
            .O(N__25398),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__4026 (
            .O(N__25395),
            .I(N__25392));
    LocalMux I__4025 (
            .O(N__25392),
            .I(N__25389));
    Span4Mux_v I__4024 (
            .O(N__25389),
            .I(N__25386));
    Odrv4 I__4023 (
            .O(N__25386),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__4022 (
            .O(N__25383),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__4021 (
            .O(N__25380),
            .I(N__25377));
    LocalMux I__4020 (
            .O(N__25377),
            .I(N__25374));
    Odrv12 I__4019 (
            .O(N__25374),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__4018 (
            .O(N__25371),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__4017 (
            .O(N__25368),
            .I(N__25365));
    LocalMux I__4016 (
            .O(N__25365),
            .I(N__25362));
    Span4Mux_v I__4015 (
            .O(N__25362),
            .I(N__25359));
    Odrv4 I__4014 (
            .O(N__25359),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__4013 (
            .O(N__25356),
            .I(bfn_8_21_0_));
    InMux I__4012 (
            .O(N__25353),
            .I(N__25350));
    LocalMux I__4011 (
            .O(N__25350),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__4010 (
            .O(N__25347),
            .I(N__25344));
    LocalMux I__4009 (
            .O(N__25344),
            .I(N__25341));
    Odrv4 I__4008 (
            .O(N__25341),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    InMux I__4007 (
            .O(N__25338),
            .I(N__25335));
    LocalMux I__4006 (
            .O(N__25335),
            .I(N__25332));
    Odrv4 I__4005 (
            .O(N__25332),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__4004 (
            .O(N__25329),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__4003 (
            .O(N__25326),
            .I(N__25323));
    LocalMux I__4002 (
            .O(N__25323),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__4001 (
            .O(N__25320),
            .I(N__25317));
    LocalMux I__4000 (
            .O(N__25317),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__3999 (
            .O(N__25314),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__3998 (
            .O(N__25311),
            .I(N__25308));
    LocalMux I__3997 (
            .O(N__25308),
            .I(N__25305));
    Span4Mux_v I__3996 (
            .O(N__25305),
            .I(N__25302));
    Odrv4 I__3995 (
            .O(N__25302),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__3994 (
            .O(N__25299),
            .I(bfn_8_20_0_));
    InMux I__3993 (
            .O(N__25296),
            .I(N__25293));
    LocalMux I__3992 (
            .O(N__25293),
            .I(N__25290));
    Odrv4 I__3991 (
            .O(N__25290),
            .I(\current_shift_inst.control_input_1_axb_18 ));
    InMux I__3990 (
            .O(N__25287),
            .I(N__25284));
    LocalMux I__3989 (
            .O(N__25284),
            .I(N__25281));
    Odrv4 I__3988 (
            .O(N__25281),
            .I(\current_shift_inst.control_input_1_axb_19 ));
    InMux I__3987 (
            .O(N__25278),
            .I(N__25275));
    LocalMux I__3986 (
            .O(N__25275),
            .I(\current_shift_inst.control_input_1_axb_24 ));
    InMux I__3985 (
            .O(N__25272),
            .I(N__25269));
    LocalMux I__3984 (
            .O(N__25269),
            .I(N__25266));
    Span4Mux_h I__3983 (
            .O(N__25266),
            .I(N__25263));
    Odrv4 I__3982 (
            .O(N__25263),
            .I(\current_shift_inst.control_input_1_axb_9 ));
    InMux I__3981 (
            .O(N__25260),
            .I(N__25257));
    LocalMux I__3980 (
            .O(N__25257),
            .I(N__25254));
    Span4Mux_v I__3979 (
            .O(N__25254),
            .I(N__25251));
    Odrv4 I__3978 (
            .O(N__25251),
            .I(\current_shift_inst.control_input_1_axb_1 ));
    InMux I__3977 (
            .O(N__25248),
            .I(N__25245));
    LocalMux I__3976 (
            .O(N__25245),
            .I(N__25242));
    Odrv4 I__3975 (
            .O(N__25242),
            .I(\current_shift_inst.control_input_1_axb_17 ));
    InMux I__3974 (
            .O(N__25239),
            .I(N__25236));
    LocalMux I__3973 (
            .O(N__25236),
            .I(N__25233));
    Span4Mux_v I__3972 (
            .O(N__25233),
            .I(N__25230));
    Odrv4 I__3971 (
            .O(N__25230),
            .I(\current_shift_inst.control_input_1_axb_4 ));
    InMux I__3970 (
            .O(N__25227),
            .I(N__25224));
    LocalMux I__3969 (
            .O(N__25224),
            .I(N__25221));
    Span4Mux_v I__3968 (
            .O(N__25221),
            .I(N__25218));
    Odrv4 I__3967 (
            .O(N__25218),
            .I(\current_shift_inst.control_input_1_axb_7 ));
    InMux I__3966 (
            .O(N__25215),
            .I(N__25212));
    LocalMux I__3965 (
            .O(N__25212),
            .I(\current_shift_inst.control_input_1_axb_16 ));
    CascadeMux I__3964 (
            .O(N__25209),
            .I(N__25206));
    InMux I__3963 (
            .O(N__25206),
            .I(N__25203));
    LocalMux I__3962 (
            .O(N__25203),
            .I(\current_shift_inst.control_input_1_axb_11 ));
    InMux I__3961 (
            .O(N__25200),
            .I(N__25197));
    LocalMux I__3960 (
            .O(N__25197),
            .I(\current_shift_inst.control_input_1_axb_8 ));
    InMux I__3959 (
            .O(N__25194),
            .I(N__25191));
    LocalMux I__3958 (
            .O(N__25191),
            .I(N__25188));
    Odrv4 I__3957 (
            .O(N__25188),
            .I(\current_shift_inst.control_input_1_axb_20 ));
    InMux I__3956 (
            .O(N__25185),
            .I(N__25182));
    LocalMux I__3955 (
            .O(N__25182),
            .I(N__25179));
    Span4Mux_h I__3954 (
            .O(N__25179),
            .I(N__25176));
    Odrv4 I__3953 (
            .O(N__25176),
            .I(\current_shift_inst.control_input_1_axb_0 ));
    InMux I__3952 (
            .O(N__25173),
            .I(N__25170));
    LocalMux I__3951 (
            .O(N__25170),
            .I(\current_shift_inst.control_input_1_axb_3 ));
    CascadeMux I__3950 (
            .O(N__25167),
            .I(N__25164));
    InMux I__3949 (
            .O(N__25164),
            .I(N__25161));
    LocalMux I__3948 (
            .O(N__25161),
            .I(N__25158));
    Odrv12 I__3947 (
            .O(N__25158),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__3946 (
            .O(N__25155),
            .I(N__25152));
    LocalMux I__3945 (
            .O(N__25152),
            .I(\current_shift_inst.control_input_1_axb_2 ));
    InMux I__3944 (
            .O(N__25149),
            .I(N__25146));
    LocalMux I__3943 (
            .O(N__25146),
            .I(\current_shift_inst.control_input_1_axb_6 ));
    InMux I__3942 (
            .O(N__25143),
            .I(N__25140));
    LocalMux I__3941 (
            .O(N__25140),
            .I(\current_shift_inst.control_input_1_axb_5 ));
    InMux I__3940 (
            .O(N__25137),
            .I(N__25134));
    LocalMux I__3939 (
            .O(N__25134),
            .I(\current_shift_inst.control_input_1_axb_14 ));
    InMux I__3938 (
            .O(N__25131),
            .I(N__25128));
    LocalMux I__3937 (
            .O(N__25128),
            .I(\current_shift_inst.control_input_1_axb_13 ));
    InMux I__3936 (
            .O(N__25125),
            .I(N__25122));
    LocalMux I__3935 (
            .O(N__25122),
            .I(\current_shift_inst.control_input_1_axb_12 ));
    InMux I__3934 (
            .O(N__25119),
            .I(N__25116));
    LocalMux I__3933 (
            .O(N__25116),
            .I(\current_shift_inst.control_input_1_axb_15 ));
    InMux I__3932 (
            .O(N__25113),
            .I(N__25110));
    LocalMux I__3931 (
            .O(N__25110),
            .I(\current_shift_inst.control_input_1_axb_10 ));
    InMux I__3930 (
            .O(N__25107),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ));
    CascadeMux I__3929 (
            .O(N__25104),
            .I(N__25101));
    InMux I__3928 (
            .O(N__25101),
            .I(N__25098));
    LocalMux I__3927 (
            .O(N__25098),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ));
    InMux I__3926 (
            .O(N__25095),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ));
    InMux I__3925 (
            .O(N__25092),
            .I(bfn_8_13_0_));
    InMux I__3924 (
            .O(N__25089),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ));
    InMux I__3923 (
            .O(N__25086),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ));
    InMux I__3922 (
            .O(N__25083),
            .I(N__25080));
    LocalMux I__3921 (
            .O(N__25080),
            .I(N__25077));
    Odrv4 I__3920 (
            .O(N__25077),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ));
    InMux I__3919 (
            .O(N__25074),
            .I(N__25071));
    LocalMux I__3918 (
            .O(N__25071),
            .I(N__25068));
    Odrv4 I__3917 (
            .O(N__25068),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ));
    InMux I__3916 (
            .O(N__25065),
            .I(N__25062));
    LocalMux I__3915 (
            .O(N__25062),
            .I(\current_shift_inst.control_input_1_axb_22 ));
    InMux I__3914 (
            .O(N__25059),
            .I(N__25056));
    LocalMux I__3913 (
            .O(N__25056),
            .I(\current_shift_inst.control_input_1_axb_21 ));
    InMux I__3912 (
            .O(N__25053),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ));
    InMux I__3911 (
            .O(N__25050),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ));
    InMux I__3910 (
            .O(N__25047),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ));
    InMux I__3909 (
            .O(N__25044),
            .I(bfn_8_12_0_));
    InMux I__3908 (
            .O(N__25041),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ));
    InMux I__3907 (
            .O(N__25038),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ));
    InMux I__3906 (
            .O(N__25035),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ));
    InMux I__3905 (
            .O(N__25032),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ));
    InMux I__3904 (
            .O(N__25029),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ));
    InMux I__3903 (
            .O(N__25026),
            .I(N__25023));
    LocalMux I__3902 (
            .O(N__25023),
            .I(N__25020));
    Odrv4 I__3901 (
            .O(N__25020),
            .I(il_min_comp2_D1));
    InMux I__3900 (
            .O(N__25017),
            .I(N__25012));
    InMux I__3899 (
            .O(N__25016),
            .I(N__25009));
    InMux I__3898 (
            .O(N__25015),
            .I(N__25006));
    LocalMux I__3897 (
            .O(N__25012),
            .I(N__25003));
    LocalMux I__3896 (
            .O(N__25009),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__3895 (
            .O(N__25006),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__3894 (
            .O(N__25003),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__3893 (
            .O(N__24996),
            .I(N__24992));
    InMux I__3892 (
            .O(N__24995),
            .I(N__24989));
    LocalMux I__3891 (
            .O(N__24992),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__3890 (
            .O(N__24989),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__3889 (
            .O(N__24984),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ));
    InMux I__3888 (
            .O(N__24981),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ));
    InMux I__3887 (
            .O(N__24978),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ));
    InMux I__3886 (
            .O(N__24975),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ));
    CascadeMux I__3885 (
            .O(N__24972),
            .I(N__24968));
    InMux I__3884 (
            .O(N__24971),
            .I(N__24965));
    InMux I__3883 (
            .O(N__24968),
            .I(N__24962));
    LocalMux I__3882 (
            .O(N__24965),
            .I(N__24959));
    LocalMux I__3881 (
            .O(N__24962),
            .I(N__24956));
    Span4Mux_h I__3880 (
            .O(N__24959),
            .I(N__24953));
    Span4Mux_h I__3879 (
            .O(N__24956),
            .I(N__24950));
    Odrv4 I__3878 (
            .O(N__24953),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    Odrv4 I__3877 (
            .O(N__24950),
            .I(\current_shift_inst.control_inputZ0Z_23 ));
    InMux I__3876 (
            .O(N__24945),
            .I(\current_shift_inst.control_input_1_cry_22 ));
    CascadeMux I__3875 (
            .O(N__24942),
            .I(N__24938));
    InMux I__3874 (
            .O(N__24941),
            .I(N__24935));
    InMux I__3873 (
            .O(N__24938),
            .I(N__24932));
    LocalMux I__3872 (
            .O(N__24935),
            .I(N__24927));
    LocalMux I__3871 (
            .O(N__24932),
            .I(N__24927));
    Odrv12 I__3870 (
            .O(N__24927),
            .I(\current_shift_inst.control_inputZ0Z_24 ));
    InMux I__3869 (
            .O(N__24924),
            .I(bfn_7_16_0_));
    InMux I__3868 (
            .O(N__24921),
            .I(\current_shift_inst.control_input_1_cry_24 ));
    CascadeMux I__3867 (
            .O(N__24918),
            .I(N__24910));
    CascadeMux I__3866 (
            .O(N__24917),
            .I(N__24906));
    CascadeMux I__3865 (
            .O(N__24916),
            .I(N__24902));
    InMux I__3864 (
            .O(N__24915),
            .I(N__24899));
    InMux I__3863 (
            .O(N__24914),
            .I(N__24884));
    InMux I__3862 (
            .O(N__24913),
            .I(N__24884));
    InMux I__3861 (
            .O(N__24910),
            .I(N__24884));
    InMux I__3860 (
            .O(N__24909),
            .I(N__24884));
    InMux I__3859 (
            .O(N__24906),
            .I(N__24884));
    InMux I__3858 (
            .O(N__24905),
            .I(N__24884));
    InMux I__3857 (
            .O(N__24902),
            .I(N__24884));
    LocalMux I__3856 (
            .O(N__24899),
            .I(N__24879));
    LocalMux I__3855 (
            .O(N__24884),
            .I(N__24879));
    Span4Mux_h I__3854 (
            .O(N__24879),
            .I(N__24876));
    Odrv4 I__3853 (
            .O(N__24876),
            .I(\current_shift_inst.control_inputZ0Z_25 ));
    CEMux I__3852 (
            .O(N__24873),
            .I(N__24868));
    CEMux I__3851 (
            .O(N__24872),
            .I(N__24863));
    CEMux I__3850 (
            .O(N__24871),
            .I(N__24858));
    LocalMux I__3849 (
            .O(N__24868),
            .I(N__24853));
    CEMux I__3848 (
            .O(N__24867),
            .I(N__24850));
    CEMux I__3847 (
            .O(N__24866),
            .I(N__24847));
    LocalMux I__3846 (
            .O(N__24863),
            .I(N__24842));
    CEMux I__3845 (
            .O(N__24862),
            .I(N__24839));
    CEMux I__3844 (
            .O(N__24861),
            .I(N__24836));
    LocalMux I__3843 (
            .O(N__24858),
            .I(N__24833));
    CEMux I__3842 (
            .O(N__24857),
            .I(N__24830));
    CEMux I__3841 (
            .O(N__24856),
            .I(N__24827));
    Span4Mux_h I__3840 (
            .O(N__24853),
            .I(N__24816));
    LocalMux I__3839 (
            .O(N__24850),
            .I(N__24816));
    LocalMux I__3838 (
            .O(N__24847),
            .I(N__24813));
    CEMux I__3837 (
            .O(N__24846),
            .I(N__24809));
    CEMux I__3836 (
            .O(N__24845),
            .I(N__24806));
    Span4Mux_v I__3835 (
            .O(N__24842),
            .I(N__24800));
    LocalMux I__3834 (
            .O(N__24839),
            .I(N__24800));
    LocalMux I__3833 (
            .O(N__24836),
            .I(N__24797));
    Span4Mux_v I__3832 (
            .O(N__24833),
            .I(N__24790));
    LocalMux I__3831 (
            .O(N__24830),
            .I(N__24790));
    LocalMux I__3830 (
            .O(N__24827),
            .I(N__24790));
    CEMux I__3829 (
            .O(N__24826),
            .I(N__24787));
    CEMux I__3828 (
            .O(N__24825),
            .I(N__24782));
    CEMux I__3827 (
            .O(N__24824),
            .I(N__24779));
    CEMux I__3826 (
            .O(N__24823),
            .I(N__24776));
    CEMux I__3825 (
            .O(N__24822),
            .I(N__24771));
    CEMux I__3824 (
            .O(N__24821),
            .I(N__24767));
    Span4Mux_v I__3823 (
            .O(N__24816),
            .I(N__24763));
    Span4Mux_h I__3822 (
            .O(N__24813),
            .I(N__24760));
    CEMux I__3821 (
            .O(N__24812),
            .I(N__24757));
    LocalMux I__3820 (
            .O(N__24809),
            .I(N__24752));
    LocalMux I__3819 (
            .O(N__24806),
            .I(N__24752));
    CEMux I__3818 (
            .O(N__24805),
            .I(N__24749));
    Span4Mux_v I__3817 (
            .O(N__24800),
            .I(N__24739));
    Span4Mux_h I__3816 (
            .O(N__24797),
            .I(N__24739));
    Span4Mux_v I__3815 (
            .O(N__24790),
            .I(N__24739));
    LocalMux I__3814 (
            .O(N__24787),
            .I(N__24739));
    CEMux I__3813 (
            .O(N__24786),
            .I(N__24736));
    CEMux I__3812 (
            .O(N__24785),
            .I(N__24733));
    LocalMux I__3811 (
            .O(N__24782),
            .I(N__24729));
    LocalMux I__3810 (
            .O(N__24779),
            .I(N__24726));
    LocalMux I__3809 (
            .O(N__24776),
            .I(N__24723));
    CEMux I__3808 (
            .O(N__24775),
            .I(N__24720));
    CEMux I__3807 (
            .O(N__24774),
            .I(N__24717));
    LocalMux I__3806 (
            .O(N__24771),
            .I(N__24713));
    CEMux I__3805 (
            .O(N__24770),
            .I(N__24710));
    LocalMux I__3804 (
            .O(N__24767),
            .I(N__24707));
    CEMux I__3803 (
            .O(N__24766),
            .I(N__24704));
    Span4Mux_v I__3802 (
            .O(N__24763),
            .I(N__24700));
    Span4Mux_v I__3801 (
            .O(N__24760),
            .I(N__24695));
    LocalMux I__3800 (
            .O(N__24757),
            .I(N__24695));
    Span4Mux_v I__3799 (
            .O(N__24752),
            .I(N__24690));
    LocalMux I__3798 (
            .O(N__24749),
            .I(N__24690));
    CEMux I__3797 (
            .O(N__24748),
            .I(N__24687));
    Span4Mux_h I__3796 (
            .O(N__24739),
            .I(N__24682));
    LocalMux I__3795 (
            .O(N__24736),
            .I(N__24682));
    LocalMux I__3794 (
            .O(N__24733),
            .I(N__24679));
    CEMux I__3793 (
            .O(N__24732),
            .I(N__24676));
    Span4Mux_v I__3792 (
            .O(N__24729),
            .I(N__24673));
    Span4Mux_h I__3791 (
            .O(N__24726),
            .I(N__24664));
    Span4Mux_v I__3790 (
            .O(N__24723),
            .I(N__24664));
    LocalMux I__3789 (
            .O(N__24720),
            .I(N__24664));
    LocalMux I__3788 (
            .O(N__24717),
            .I(N__24664));
    CEMux I__3787 (
            .O(N__24716),
            .I(N__24661));
    Span4Mux_h I__3786 (
            .O(N__24713),
            .I(N__24652));
    LocalMux I__3785 (
            .O(N__24710),
            .I(N__24652));
    Span4Mux_v I__3784 (
            .O(N__24707),
            .I(N__24652));
    LocalMux I__3783 (
            .O(N__24704),
            .I(N__24652));
    CEMux I__3782 (
            .O(N__24703),
            .I(N__24649));
    Span4Mux_v I__3781 (
            .O(N__24700),
            .I(N__24646));
    Span4Mux_h I__3780 (
            .O(N__24695),
            .I(N__24643));
    Span4Mux_v I__3779 (
            .O(N__24690),
            .I(N__24640));
    LocalMux I__3778 (
            .O(N__24687),
            .I(N__24637));
    Span4Mux_v I__3777 (
            .O(N__24682),
            .I(N__24634));
    Span4Mux_v I__3776 (
            .O(N__24679),
            .I(N__24629));
    LocalMux I__3775 (
            .O(N__24676),
            .I(N__24629));
    Span4Mux_h I__3774 (
            .O(N__24673),
            .I(N__24622));
    Span4Mux_v I__3773 (
            .O(N__24664),
            .I(N__24622));
    LocalMux I__3772 (
            .O(N__24661),
            .I(N__24622));
    Span4Mux_v I__3771 (
            .O(N__24652),
            .I(N__24617));
    LocalMux I__3770 (
            .O(N__24649),
            .I(N__24617));
    Span4Mux_h I__3769 (
            .O(N__24646),
            .I(N__24614));
    Span4Mux_v I__3768 (
            .O(N__24643),
            .I(N__24609));
    Span4Mux_h I__3767 (
            .O(N__24640),
            .I(N__24609));
    Span4Mux_h I__3766 (
            .O(N__24637),
            .I(N__24606));
    Span4Mux_s2_h I__3765 (
            .O(N__24634),
            .I(N__24601));
    Span4Mux_v I__3764 (
            .O(N__24629),
            .I(N__24601));
    Span4Mux_v I__3763 (
            .O(N__24622),
            .I(N__24596));
    Span4Mux_h I__3762 (
            .O(N__24617),
            .I(N__24596));
    Odrv4 I__3761 (
            .O(N__24614),
            .I(N_748_g));
    Odrv4 I__3760 (
            .O(N__24609),
            .I(N_748_g));
    Odrv4 I__3759 (
            .O(N__24606),
            .I(N_748_g));
    Odrv4 I__3758 (
            .O(N__24601),
            .I(N_748_g));
    Odrv4 I__3757 (
            .O(N__24596),
            .I(N_748_g));
    InMux I__3756 (
            .O(N__24585),
            .I(N__24582));
    LocalMux I__3755 (
            .O(N__24582),
            .I(N__24579));
    Sp12to4 I__3754 (
            .O(N__24579),
            .I(N__24576));
    Odrv12 I__3753 (
            .O(N__24576),
            .I(\current_shift_inst.control_input_1_axb_23 ));
    InMux I__3752 (
            .O(N__24573),
            .I(N__24570));
    LocalMux I__3751 (
            .O(N__24570),
            .I(N__24567));
    Odrv12 I__3750 (
            .O(N__24567),
            .I(il_max_comp1_c));
    InMux I__3749 (
            .O(N__24564),
            .I(N__24561));
    LocalMux I__3748 (
            .O(N__24561),
            .I(N__24558));
    Span4Mux_h I__3747 (
            .O(N__24558),
            .I(N__24555));
    Span4Mux_v I__3746 (
            .O(N__24555),
            .I(N__24552));
    Odrv4 I__3745 (
            .O(N__24552),
            .I(il_min_comp2_c));
    InMux I__3744 (
            .O(N__24549),
            .I(N__24545));
    InMux I__3743 (
            .O(N__24548),
            .I(N__24542));
    LocalMux I__3742 (
            .O(N__24545),
            .I(N__24537));
    LocalMux I__3741 (
            .O(N__24542),
            .I(N__24537));
    Span4Mux_h I__3740 (
            .O(N__24537),
            .I(N__24534));
    Odrv4 I__3739 (
            .O(N__24534),
            .I(\current_shift_inst.control_inputZ0Z_15 ));
    InMux I__3738 (
            .O(N__24531),
            .I(\current_shift_inst.control_input_1_cry_14 ));
    CascadeMux I__3737 (
            .O(N__24528),
            .I(N__24524));
    InMux I__3736 (
            .O(N__24527),
            .I(N__24521));
    InMux I__3735 (
            .O(N__24524),
            .I(N__24518));
    LocalMux I__3734 (
            .O(N__24521),
            .I(N__24515));
    LocalMux I__3733 (
            .O(N__24518),
            .I(N__24512));
    Span4Mux_h I__3732 (
            .O(N__24515),
            .I(N__24509));
    Span4Mux_h I__3731 (
            .O(N__24512),
            .I(N__24506));
    Odrv4 I__3730 (
            .O(N__24509),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    Odrv4 I__3729 (
            .O(N__24506),
            .I(\current_shift_inst.control_inputZ0Z_16 ));
    InMux I__3728 (
            .O(N__24501),
            .I(bfn_7_15_0_));
    CascadeMux I__3727 (
            .O(N__24498),
            .I(N__24494));
    InMux I__3726 (
            .O(N__24497),
            .I(N__24491));
    InMux I__3725 (
            .O(N__24494),
            .I(N__24488));
    LocalMux I__3724 (
            .O(N__24491),
            .I(N__24483));
    LocalMux I__3723 (
            .O(N__24488),
            .I(N__24483));
    Odrv12 I__3722 (
            .O(N__24483),
            .I(\current_shift_inst.control_inputZ0Z_17 ));
    InMux I__3721 (
            .O(N__24480),
            .I(\current_shift_inst.control_input_1_cry_16 ));
    CascadeMux I__3720 (
            .O(N__24477),
            .I(N__24473));
    InMux I__3719 (
            .O(N__24476),
            .I(N__24470));
    InMux I__3718 (
            .O(N__24473),
            .I(N__24467));
    LocalMux I__3717 (
            .O(N__24470),
            .I(N__24464));
    LocalMux I__3716 (
            .O(N__24467),
            .I(N__24461));
    Odrv12 I__3715 (
            .O(N__24464),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    Odrv4 I__3714 (
            .O(N__24461),
            .I(\current_shift_inst.control_inputZ0Z_18 ));
    InMux I__3713 (
            .O(N__24456),
            .I(\current_shift_inst.control_input_1_cry_17 ));
    CascadeMux I__3712 (
            .O(N__24453),
            .I(N__24449));
    InMux I__3711 (
            .O(N__24452),
            .I(N__24446));
    InMux I__3710 (
            .O(N__24449),
            .I(N__24443));
    LocalMux I__3709 (
            .O(N__24446),
            .I(N__24438));
    LocalMux I__3708 (
            .O(N__24443),
            .I(N__24438));
    Odrv12 I__3707 (
            .O(N__24438),
            .I(\current_shift_inst.control_inputZ0Z_19 ));
    InMux I__3706 (
            .O(N__24435),
            .I(\current_shift_inst.control_input_1_cry_18 ));
    CascadeMux I__3705 (
            .O(N__24432),
            .I(N__24428));
    InMux I__3704 (
            .O(N__24431),
            .I(N__24425));
    InMux I__3703 (
            .O(N__24428),
            .I(N__24422));
    LocalMux I__3702 (
            .O(N__24425),
            .I(N__24419));
    LocalMux I__3701 (
            .O(N__24422),
            .I(N__24416));
    Odrv12 I__3700 (
            .O(N__24419),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    Odrv4 I__3699 (
            .O(N__24416),
            .I(\current_shift_inst.control_inputZ0Z_20 ));
    InMux I__3698 (
            .O(N__24411),
            .I(\current_shift_inst.control_input_1_cry_19 ));
    InMux I__3697 (
            .O(N__24408),
            .I(N__24404));
    CascadeMux I__3696 (
            .O(N__24407),
            .I(N__24401));
    LocalMux I__3695 (
            .O(N__24404),
            .I(N__24398));
    InMux I__3694 (
            .O(N__24401),
            .I(N__24395));
    Span4Mux_v I__3693 (
            .O(N__24398),
            .I(N__24390));
    LocalMux I__3692 (
            .O(N__24395),
            .I(N__24390));
    Odrv4 I__3691 (
            .O(N__24390),
            .I(\current_shift_inst.control_inputZ0Z_21 ));
    InMux I__3690 (
            .O(N__24387),
            .I(\current_shift_inst.control_input_1_cry_20 ));
    CascadeMux I__3689 (
            .O(N__24384),
            .I(N__24380));
    InMux I__3688 (
            .O(N__24383),
            .I(N__24377));
    InMux I__3687 (
            .O(N__24380),
            .I(N__24374));
    LocalMux I__3686 (
            .O(N__24377),
            .I(N__24369));
    LocalMux I__3685 (
            .O(N__24374),
            .I(N__24369));
    Odrv12 I__3684 (
            .O(N__24369),
            .I(\current_shift_inst.control_inputZ0Z_22 ));
    InMux I__3683 (
            .O(N__24366),
            .I(\current_shift_inst.control_input_1_cry_21 ));
    CascadeMux I__3682 (
            .O(N__24363),
            .I(N__24359));
    InMux I__3681 (
            .O(N__24362),
            .I(N__24356));
    InMux I__3680 (
            .O(N__24359),
            .I(N__24353));
    LocalMux I__3679 (
            .O(N__24356),
            .I(N__24348));
    LocalMux I__3678 (
            .O(N__24353),
            .I(N__24348));
    Span4Mux_h I__3677 (
            .O(N__24348),
            .I(N__24345));
    Odrv4 I__3676 (
            .O(N__24345),
            .I(\current_shift_inst.control_inputZ0Z_6 ));
    InMux I__3675 (
            .O(N__24342),
            .I(\current_shift_inst.control_input_1_cry_5 ));
    CascadeMux I__3674 (
            .O(N__24339),
            .I(N__24335));
    InMux I__3673 (
            .O(N__24338),
            .I(N__24332));
    InMux I__3672 (
            .O(N__24335),
            .I(N__24329));
    LocalMux I__3671 (
            .O(N__24332),
            .I(N__24324));
    LocalMux I__3670 (
            .O(N__24329),
            .I(N__24324));
    Span4Mux_h I__3669 (
            .O(N__24324),
            .I(N__24321));
    Odrv4 I__3668 (
            .O(N__24321),
            .I(\current_shift_inst.control_inputZ0Z_7 ));
    InMux I__3667 (
            .O(N__24318),
            .I(\current_shift_inst.control_input_1_cry_6 ));
    CascadeMux I__3666 (
            .O(N__24315),
            .I(N__24311));
    InMux I__3665 (
            .O(N__24314),
            .I(N__24308));
    InMux I__3664 (
            .O(N__24311),
            .I(N__24305));
    LocalMux I__3663 (
            .O(N__24308),
            .I(N__24300));
    LocalMux I__3662 (
            .O(N__24305),
            .I(N__24300));
    Span4Mux_h I__3661 (
            .O(N__24300),
            .I(N__24297));
    Odrv4 I__3660 (
            .O(N__24297),
            .I(\current_shift_inst.control_inputZ0Z_8 ));
    InMux I__3659 (
            .O(N__24294),
            .I(bfn_7_14_0_));
    CascadeMux I__3658 (
            .O(N__24291),
            .I(N__24287));
    InMux I__3657 (
            .O(N__24290),
            .I(N__24284));
    InMux I__3656 (
            .O(N__24287),
            .I(N__24281));
    LocalMux I__3655 (
            .O(N__24284),
            .I(N__24276));
    LocalMux I__3654 (
            .O(N__24281),
            .I(N__24276));
    Span4Mux_h I__3653 (
            .O(N__24276),
            .I(N__24273));
    Odrv4 I__3652 (
            .O(N__24273),
            .I(\current_shift_inst.control_inputZ0Z_9 ));
    InMux I__3651 (
            .O(N__24270),
            .I(\current_shift_inst.control_input_1_cry_8 ));
    InMux I__3650 (
            .O(N__24267),
            .I(N__24263));
    CascadeMux I__3649 (
            .O(N__24266),
            .I(N__24260));
    LocalMux I__3648 (
            .O(N__24263),
            .I(N__24257));
    InMux I__3647 (
            .O(N__24260),
            .I(N__24254));
    Span4Mux_v I__3646 (
            .O(N__24257),
            .I(N__24249));
    LocalMux I__3645 (
            .O(N__24254),
            .I(N__24249));
    Odrv4 I__3644 (
            .O(N__24249),
            .I(\current_shift_inst.control_inputZ0Z_10 ));
    InMux I__3643 (
            .O(N__24246),
            .I(\current_shift_inst.control_input_1_cry_9 ));
    InMux I__3642 (
            .O(N__24243),
            .I(N__24239));
    InMux I__3641 (
            .O(N__24242),
            .I(N__24236));
    LocalMux I__3640 (
            .O(N__24239),
            .I(N__24231));
    LocalMux I__3639 (
            .O(N__24236),
            .I(N__24231));
    Span4Mux_h I__3638 (
            .O(N__24231),
            .I(N__24228));
    Odrv4 I__3637 (
            .O(N__24228),
            .I(\current_shift_inst.control_inputZ0Z_11 ));
    InMux I__3636 (
            .O(N__24225),
            .I(\current_shift_inst.control_input_1_cry_10 ));
    CascadeMux I__3635 (
            .O(N__24222),
            .I(N__24218));
    InMux I__3634 (
            .O(N__24221),
            .I(N__24215));
    InMux I__3633 (
            .O(N__24218),
            .I(N__24212));
    LocalMux I__3632 (
            .O(N__24215),
            .I(N__24209));
    LocalMux I__3631 (
            .O(N__24212),
            .I(N__24206));
    Odrv12 I__3630 (
            .O(N__24209),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    Odrv4 I__3629 (
            .O(N__24206),
            .I(\current_shift_inst.control_inputZ0Z_12 ));
    InMux I__3628 (
            .O(N__24201),
            .I(\current_shift_inst.control_input_1_cry_11 ));
    InMux I__3627 (
            .O(N__24198),
            .I(N__24194));
    CascadeMux I__3626 (
            .O(N__24197),
            .I(N__24191));
    LocalMux I__3625 (
            .O(N__24194),
            .I(N__24188));
    InMux I__3624 (
            .O(N__24191),
            .I(N__24185));
    Span4Mux_v I__3623 (
            .O(N__24188),
            .I(N__24180));
    LocalMux I__3622 (
            .O(N__24185),
            .I(N__24180));
    Odrv4 I__3621 (
            .O(N__24180),
            .I(\current_shift_inst.control_inputZ0Z_13 ));
    InMux I__3620 (
            .O(N__24177),
            .I(\current_shift_inst.control_input_1_cry_12 ));
    CascadeMux I__3619 (
            .O(N__24174),
            .I(N__24170));
    InMux I__3618 (
            .O(N__24173),
            .I(N__24167));
    InMux I__3617 (
            .O(N__24170),
            .I(N__24164));
    LocalMux I__3616 (
            .O(N__24167),
            .I(N__24159));
    LocalMux I__3615 (
            .O(N__24164),
            .I(N__24159));
    Odrv12 I__3614 (
            .O(N__24159),
            .I(\current_shift_inst.control_inputZ0Z_14 ));
    InMux I__3613 (
            .O(N__24156),
            .I(\current_shift_inst.control_input_1_cry_13 ));
    CascadeMux I__3612 (
            .O(N__24153),
            .I(\phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa_cascade_ ));
    CascadeMux I__3611 (
            .O(N__24150),
            .I(N__24147));
    InMux I__3610 (
            .O(N__24147),
            .I(N__24144));
    LocalMux I__3609 (
            .O(N__24144),
            .I(N__24141));
    Span4Mux_s3_h I__3608 (
            .O(N__24141),
            .I(N__24138));
    Span4Mux_h I__3607 (
            .O(N__24138),
            .I(N__24135));
    Odrv4 I__3606 (
            .O(N__24135),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__3605 (
            .O(N__24132),
            .I(N__24128));
    CascadeMux I__3604 (
            .O(N__24131),
            .I(N__24124));
    LocalMux I__3603 (
            .O(N__24128),
            .I(N__24121));
    InMux I__3602 (
            .O(N__24127),
            .I(N__24118));
    InMux I__3601 (
            .O(N__24124),
            .I(N__24115));
    Span4Mux_v I__3600 (
            .O(N__24121),
            .I(N__24112));
    LocalMux I__3599 (
            .O(N__24118),
            .I(N__24107));
    LocalMux I__3598 (
            .O(N__24115),
            .I(N__24107));
    Span4Mux_h I__3597 (
            .O(N__24112),
            .I(N__24104));
    Span4Mux_h I__3596 (
            .O(N__24107),
            .I(N__24101));
    Odrv4 I__3595 (
            .O(N__24104),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    Odrv4 I__3594 (
            .O(N__24101),
            .I(\current_shift_inst.control_inputZ0Z_0 ));
    CascadeMux I__3593 (
            .O(N__24096),
            .I(N__24092));
    InMux I__3592 (
            .O(N__24095),
            .I(N__24089));
    InMux I__3591 (
            .O(N__24092),
            .I(N__24086));
    LocalMux I__3590 (
            .O(N__24089),
            .I(N__24081));
    LocalMux I__3589 (
            .O(N__24086),
            .I(N__24081));
    Span4Mux_h I__3588 (
            .O(N__24081),
            .I(N__24078));
    Odrv4 I__3587 (
            .O(N__24078),
            .I(\current_shift_inst.control_inputZ0Z_1 ));
    InMux I__3586 (
            .O(N__24075),
            .I(\current_shift_inst.control_input_1_cry_0 ));
    CascadeMux I__3585 (
            .O(N__24072),
            .I(N__24069));
    InMux I__3584 (
            .O(N__24069),
            .I(N__24065));
    InMux I__3583 (
            .O(N__24068),
            .I(N__24062));
    LocalMux I__3582 (
            .O(N__24065),
            .I(N__24059));
    LocalMux I__3581 (
            .O(N__24062),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    Odrv12 I__3580 (
            .O(N__24059),
            .I(\current_shift_inst.control_inputZ0Z_2 ));
    InMux I__3579 (
            .O(N__24054),
            .I(\current_shift_inst.control_input_1_cry_1 ));
    CascadeMux I__3578 (
            .O(N__24051),
            .I(N__24047));
    InMux I__3577 (
            .O(N__24050),
            .I(N__24044));
    InMux I__3576 (
            .O(N__24047),
            .I(N__24041));
    LocalMux I__3575 (
            .O(N__24044),
            .I(N__24036));
    LocalMux I__3574 (
            .O(N__24041),
            .I(N__24036));
    Odrv12 I__3573 (
            .O(N__24036),
            .I(\current_shift_inst.control_inputZ0Z_3 ));
    InMux I__3572 (
            .O(N__24033),
            .I(\current_shift_inst.control_input_1_cry_2 ));
    CascadeMux I__3571 (
            .O(N__24030),
            .I(N__24026));
    InMux I__3570 (
            .O(N__24029),
            .I(N__24023));
    InMux I__3569 (
            .O(N__24026),
            .I(N__24020));
    LocalMux I__3568 (
            .O(N__24023),
            .I(N__24015));
    LocalMux I__3567 (
            .O(N__24020),
            .I(N__24015));
    Odrv12 I__3566 (
            .O(N__24015),
            .I(\current_shift_inst.control_inputZ0Z_4 ));
    InMux I__3565 (
            .O(N__24012),
            .I(\current_shift_inst.control_input_1_cry_3 ));
    CascadeMux I__3564 (
            .O(N__24009),
            .I(N__24005));
    InMux I__3563 (
            .O(N__24008),
            .I(N__24002));
    InMux I__3562 (
            .O(N__24005),
            .I(N__23999));
    LocalMux I__3561 (
            .O(N__24002),
            .I(N__23996));
    LocalMux I__3560 (
            .O(N__23999),
            .I(N__23993));
    Odrv12 I__3559 (
            .O(N__23996),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    Odrv4 I__3558 (
            .O(N__23993),
            .I(\current_shift_inst.control_inputZ0Z_5 ));
    InMux I__3557 (
            .O(N__23988),
            .I(\current_shift_inst.control_input_1_cry_4 ));
    CascadeMux I__3556 (
            .O(N__23985),
            .I(N__23982));
    InMux I__3555 (
            .O(N__23982),
            .I(N__23979));
    LocalMux I__3554 (
            .O(N__23979),
            .I(N__23975));
    InMux I__3553 (
            .O(N__23978),
            .I(N__23970));
    Span4Mux_v I__3552 (
            .O(N__23975),
            .I(N__23967));
    InMux I__3551 (
            .O(N__23974),
            .I(N__23964));
    CascadeMux I__3550 (
            .O(N__23973),
            .I(N__23961));
    LocalMux I__3549 (
            .O(N__23970),
            .I(N__23958));
    Span4Mux_h I__3548 (
            .O(N__23967),
            .I(N__23953));
    LocalMux I__3547 (
            .O(N__23964),
            .I(N__23953));
    InMux I__3546 (
            .O(N__23961),
            .I(N__23950));
    Odrv4 I__3545 (
            .O(N__23958),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__3544 (
            .O(N__23953),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3543 (
            .O(N__23950),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__3542 (
            .O(N__23943),
            .I(N__23940));
    InMux I__3541 (
            .O(N__23940),
            .I(N__23937));
    LocalMux I__3540 (
            .O(N__23937),
            .I(N__23934));
    Span4Mux_h I__3539 (
            .O(N__23934),
            .I(N__23931));
    Odrv4 I__3538 (
            .O(N__23931),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__3537 (
            .O(N__23928),
            .I(N__23925));
    LocalMux I__3536 (
            .O(N__23925),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__3535 (
            .O(N__23922),
            .I(N__23911));
    CascadeMux I__3534 (
            .O(N__23921),
            .I(N__23908));
    CascadeMux I__3533 (
            .O(N__23920),
            .I(N__23902));
    InMux I__3532 (
            .O(N__23919),
            .I(N__23892));
    InMux I__3531 (
            .O(N__23918),
            .I(N__23892));
    InMux I__3530 (
            .O(N__23917),
            .I(N__23889));
    InMux I__3529 (
            .O(N__23916),
            .I(N__23882));
    InMux I__3528 (
            .O(N__23915),
            .I(N__23882));
    InMux I__3527 (
            .O(N__23914),
            .I(N__23882));
    InMux I__3526 (
            .O(N__23911),
            .I(N__23871));
    InMux I__3525 (
            .O(N__23908),
            .I(N__23871));
    InMux I__3524 (
            .O(N__23907),
            .I(N__23871));
    InMux I__3523 (
            .O(N__23906),
            .I(N__23871));
    InMux I__3522 (
            .O(N__23905),
            .I(N__23871));
    InMux I__3521 (
            .O(N__23902),
            .I(N__23855));
    InMux I__3520 (
            .O(N__23901),
            .I(N__23855));
    InMux I__3519 (
            .O(N__23900),
            .I(N__23855));
    CascadeMux I__3518 (
            .O(N__23899),
            .I(N__23852));
    CascadeMux I__3517 (
            .O(N__23898),
            .I(N__23848));
    CascadeMux I__3516 (
            .O(N__23897),
            .I(N__23845));
    LocalMux I__3515 (
            .O(N__23892),
            .I(N__23834));
    LocalMux I__3514 (
            .O(N__23889),
            .I(N__23834));
    LocalMux I__3513 (
            .O(N__23882),
            .I(N__23834));
    LocalMux I__3512 (
            .O(N__23871),
            .I(N__23834));
    InMux I__3511 (
            .O(N__23870),
            .I(N__23827));
    InMux I__3510 (
            .O(N__23869),
            .I(N__23827));
    InMux I__3509 (
            .O(N__23868),
            .I(N__23827));
    InMux I__3508 (
            .O(N__23867),
            .I(N__23818));
    InMux I__3507 (
            .O(N__23866),
            .I(N__23818));
    InMux I__3506 (
            .O(N__23865),
            .I(N__23818));
    InMux I__3505 (
            .O(N__23864),
            .I(N__23818));
    InMux I__3504 (
            .O(N__23863),
            .I(N__23815));
    InMux I__3503 (
            .O(N__23862),
            .I(N__23812));
    LocalMux I__3502 (
            .O(N__23855),
            .I(N__23809));
    InMux I__3501 (
            .O(N__23852),
            .I(N__23796));
    InMux I__3500 (
            .O(N__23851),
            .I(N__23796));
    InMux I__3499 (
            .O(N__23848),
            .I(N__23796));
    InMux I__3498 (
            .O(N__23845),
            .I(N__23796));
    InMux I__3497 (
            .O(N__23844),
            .I(N__23796));
    InMux I__3496 (
            .O(N__23843),
            .I(N__23796));
    Span4Mux_v I__3495 (
            .O(N__23834),
            .I(N__23785));
    LocalMux I__3494 (
            .O(N__23827),
            .I(N__23785));
    LocalMux I__3493 (
            .O(N__23818),
            .I(N__23785));
    LocalMux I__3492 (
            .O(N__23815),
            .I(N__23785));
    LocalMux I__3491 (
            .O(N__23812),
            .I(N__23782));
    Span4Mux_v I__3490 (
            .O(N__23809),
            .I(N__23777));
    LocalMux I__3489 (
            .O(N__23796),
            .I(N__23777));
    InMux I__3488 (
            .O(N__23795),
            .I(N__23774));
    InMux I__3487 (
            .O(N__23794),
            .I(N__23771));
    Odrv4 I__3486 (
            .O(N__23785),
            .I(\current_shift_inst.PI_CTRL.N_170 ));
    Odrv4 I__3485 (
            .O(N__23782),
            .I(\current_shift_inst.PI_CTRL.N_170 ));
    Odrv4 I__3484 (
            .O(N__23777),
            .I(\current_shift_inst.PI_CTRL.N_170 ));
    LocalMux I__3483 (
            .O(N__23774),
            .I(\current_shift_inst.PI_CTRL.N_170 ));
    LocalMux I__3482 (
            .O(N__23771),
            .I(\current_shift_inst.PI_CTRL.N_170 ));
    InMux I__3481 (
            .O(N__23760),
            .I(N__23748));
    InMux I__3480 (
            .O(N__23759),
            .I(N__23748));
    InMux I__3479 (
            .O(N__23758),
            .I(N__23748));
    InMux I__3478 (
            .O(N__23757),
            .I(N__23742));
    InMux I__3477 (
            .O(N__23756),
            .I(N__23737));
    InMux I__3476 (
            .O(N__23755),
            .I(N__23737));
    LocalMux I__3475 (
            .O(N__23748),
            .I(N__23725));
    InMux I__3474 (
            .O(N__23747),
            .I(N__23720));
    InMux I__3473 (
            .O(N__23746),
            .I(N__23720));
    InMux I__3472 (
            .O(N__23745),
            .I(N__23717));
    LocalMux I__3471 (
            .O(N__23742),
            .I(N__23714));
    LocalMux I__3470 (
            .O(N__23737),
            .I(N__23711));
    InMux I__3469 (
            .O(N__23736),
            .I(N__23702));
    InMux I__3468 (
            .O(N__23735),
            .I(N__23702));
    InMux I__3467 (
            .O(N__23734),
            .I(N__23702));
    InMux I__3466 (
            .O(N__23733),
            .I(N__23702));
    InMux I__3465 (
            .O(N__23732),
            .I(N__23691));
    InMux I__3464 (
            .O(N__23731),
            .I(N__23691));
    InMux I__3463 (
            .O(N__23730),
            .I(N__23691));
    InMux I__3462 (
            .O(N__23729),
            .I(N__23691));
    InMux I__3461 (
            .O(N__23728),
            .I(N__23691));
    Span4Mux_h I__3460 (
            .O(N__23725),
            .I(N__23675));
    LocalMux I__3459 (
            .O(N__23720),
            .I(N__23670));
    LocalMux I__3458 (
            .O(N__23717),
            .I(N__23670));
    Span4Mux_v I__3457 (
            .O(N__23714),
            .I(N__23661));
    Span4Mux_v I__3456 (
            .O(N__23711),
            .I(N__23661));
    LocalMux I__3455 (
            .O(N__23702),
            .I(N__23661));
    LocalMux I__3454 (
            .O(N__23691),
            .I(N__23661));
    InMux I__3453 (
            .O(N__23690),
            .I(N__23648));
    InMux I__3452 (
            .O(N__23689),
            .I(N__23648));
    InMux I__3451 (
            .O(N__23688),
            .I(N__23648));
    InMux I__3450 (
            .O(N__23687),
            .I(N__23648));
    InMux I__3449 (
            .O(N__23686),
            .I(N__23648));
    InMux I__3448 (
            .O(N__23685),
            .I(N__23648));
    InMux I__3447 (
            .O(N__23684),
            .I(N__23633));
    InMux I__3446 (
            .O(N__23683),
            .I(N__23633));
    InMux I__3445 (
            .O(N__23682),
            .I(N__23633));
    InMux I__3444 (
            .O(N__23681),
            .I(N__23633));
    InMux I__3443 (
            .O(N__23680),
            .I(N__23633));
    InMux I__3442 (
            .O(N__23679),
            .I(N__23633));
    InMux I__3441 (
            .O(N__23678),
            .I(N__23633));
    Odrv4 I__3440 (
            .O(N__23675),
            .I(\current_shift_inst.PI_CTRL.N_171 ));
    Odrv4 I__3439 (
            .O(N__23670),
            .I(\current_shift_inst.PI_CTRL.N_171 ));
    Odrv4 I__3438 (
            .O(N__23661),
            .I(\current_shift_inst.PI_CTRL.N_171 ));
    LocalMux I__3437 (
            .O(N__23648),
            .I(\current_shift_inst.PI_CTRL.N_171 ));
    LocalMux I__3436 (
            .O(N__23633),
            .I(\current_shift_inst.PI_CTRL.N_171 ));
    CascadeMux I__3435 (
            .O(N__23622),
            .I(N__23614));
    CascadeMux I__3434 (
            .O(N__23621),
            .I(N__23607));
    CascadeMux I__3433 (
            .O(N__23620),
            .I(N__23604));
    CascadeMux I__3432 (
            .O(N__23619),
            .I(N__23596));
    CascadeMux I__3431 (
            .O(N__23618),
            .I(N__23593));
    CascadeMux I__3430 (
            .O(N__23617),
            .I(N__23590));
    InMux I__3429 (
            .O(N__23614),
            .I(N__23585));
    CascadeMux I__3428 (
            .O(N__23613),
            .I(N__23576));
    CascadeMux I__3427 (
            .O(N__23612),
            .I(N__23573));
    CascadeMux I__3426 (
            .O(N__23611),
            .I(N__23570));
    CascadeMux I__3425 (
            .O(N__23610),
            .I(N__23567));
    InMux I__3424 (
            .O(N__23607),
            .I(N__23558));
    InMux I__3423 (
            .O(N__23604),
            .I(N__23558));
    InMux I__3422 (
            .O(N__23603),
            .I(N__23558));
    CascadeMux I__3421 (
            .O(N__23602),
            .I(N__23554));
    CascadeMux I__3420 (
            .O(N__23601),
            .I(N__23551));
    CascadeMux I__3419 (
            .O(N__23600),
            .I(N__23548));
    CascadeMux I__3418 (
            .O(N__23599),
            .I(N__23545));
    InMux I__3417 (
            .O(N__23596),
            .I(N__23539));
    InMux I__3416 (
            .O(N__23593),
            .I(N__23532));
    InMux I__3415 (
            .O(N__23590),
            .I(N__23532));
    InMux I__3414 (
            .O(N__23589),
            .I(N__23532));
    InMux I__3413 (
            .O(N__23588),
            .I(N__23529));
    LocalMux I__3412 (
            .O(N__23585),
            .I(N__23526));
    CascadeMux I__3411 (
            .O(N__23584),
            .I(N__23521));
    CascadeMux I__3410 (
            .O(N__23583),
            .I(N__23518));
    CascadeMux I__3409 (
            .O(N__23582),
            .I(N__23515));
    CascadeMux I__3408 (
            .O(N__23581),
            .I(N__23512));
    CascadeMux I__3407 (
            .O(N__23580),
            .I(N__23509));
    InMux I__3406 (
            .O(N__23579),
            .I(N__23505));
    InMux I__3405 (
            .O(N__23576),
            .I(N__23502));
    InMux I__3404 (
            .O(N__23573),
            .I(N__23491));
    InMux I__3403 (
            .O(N__23570),
            .I(N__23491));
    InMux I__3402 (
            .O(N__23567),
            .I(N__23491));
    InMux I__3401 (
            .O(N__23566),
            .I(N__23491));
    InMux I__3400 (
            .O(N__23565),
            .I(N__23491));
    LocalMux I__3399 (
            .O(N__23558),
            .I(N__23488));
    CascadeMux I__3398 (
            .O(N__23557),
            .I(N__23485));
    InMux I__3397 (
            .O(N__23554),
            .I(N__23472));
    InMux I__3396 (
            .O(N__23551),
            .I(N__23472));
    InMux I__3395 (
            .O(N__23548),
            .I(N__23472));
    InMux I__3394 (
            .O(N__23545),
            .I(N__23472));
    InMux I__3393 (
            .O(N__23544),
            .I(N__23472));
    InMux I__3392 (
            .O(N__23543),
            .I(N__23472));
    InMux I__3391 (
            .O(N__23542),
            .I(N__23469));
    LocalMux I__3390 (
            .O(N__23539),
            .I(N__23460));
    LocalMux I__3389 (
            .O(N__23532),
            .I(N__23460));
    LocalMux I__3388 (
            .O(N__23529),
            .I(N__23460));
    Span4Mux_h I__3387 (
            .O(N__23526),
            .I(N__23460));
    InMux I__3386 (
            .O(N__23525),
            .I(N__23457));
    CascadeMux I__3385 (
            .O(N__23524),
            .I(N__23454));
    InMux I__3384 (
            .O(N__23521),
            .I(N__23449));
    InMux I__3383 (
            .O(N__23518),
            .I(N__23449));
    InMux I__3382 (
            .O(N__23515),
            .I(N__23440));
    InMux I__3381 (
            .O(N__23512),
            .I(N__23440));
    InMux I__3380 (
            .O(N__23509),
            .I(N__23440));
    InMux I__3379 (
            .O(N__23508),
            .I(N__23440));
    LocalMux I__3378 (
            .O(N__23505),
            .I(N__23437));
    LocalMux I__3377 (
            .O(N__23502),
            .I(N__23432));
    LocalMux I__3376 (
            .O(N__23491),
            .I(N__23432));
    Span4Mux_h I__3375 (
            .O(N__23488),
            .I(N__23429));
    InMux I__3374 (
            .O(N__23485),
            .I(N__23426));
    LocalMux I__3373 (
            .O(N__23472),
            .I(N__23417));
    LocalMux I__3372 (
            .O(N__23469),
            .I(N__23417));
    Sp12to4 I__3371 (
            .O(N__23460),
            .I(N__23417));
    LocalMux I__3370 (
            .O(N__23457),
            .I(N__23417));
    InMux I__3369 (
            .O(N__23454),
            .I(N__23414));
    LocalMux I__3368 (
            .O(N__23449),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3367 (
            .O(N__23440),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3366 (
            .O(N__23437),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3365 (
            .O(N__23432),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3364 (
            .O(N__23429),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3363 (
            .O(N__23426),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3362 (
            .O(N__23417),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3361 (
            .O(N__23414),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__3360 (
            .O(N__23397),
            .I(N__23394));
    LocalMux I__3359 (
            .O(N__23394),
            .I(N__23391));
    Span4Mux_h I__3358 (
            .O(N__23391),
            .I(N__23388));
    Odrv4 I__3357 (
            .O(N__23388),
            .I(il_max_comp2_c));
    InMux I__3356 (
            .O(N__23385),
            .I(N__23382));
    LocalMux I__3355 (
            .O(N__23382),
            .I(N__23377));
    InMux I__3354 (
            .O(N__23381),
            .I(N__23374));
    InMux I__3353 (
            .O(N__23380),
            .I(N__23371));
    Span4Mux_v I__3352 (
            .O(N__23377),
            .I(N__23368));
    LocalMux I__3351 (
            .O(N__23374),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__3350 (
            .O(N__23371),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__3349 (
            .O(N__23368),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__3348 (
            .O(N__23361),
            .I(N__23358));
    LocalMux I__3347 (
            .O(N__23358),
            .I(N__23353));
    InMux I__3346 (
            .O(N__23357),
            .I(N__23350));
    InMux I__3345 (
            .O(N__23356),
            .I(N__23347));
    Span4Mux_v I__3344 (
            .O(N__23353),
            .I(N__23344));
    LocalMux I__3343 (
            .O(N__23350),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__3342 (
            .O(N__23347),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__3341 (
            .O(N__23344),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__3340 (
            .O(N__23337),
            .I(N__23333));
    InMux I__3339 (
            .O(N__23336),
            .I(N__23329));
    LocalMux I__3338 (
            .O(N__23333),
            .I(N__23326));
    InMux I__3337 (
            .O(N__23332),
            .I(N__23323));
    LocalMux I__3336 (
            .O(N__23329),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__3335 (
            .O(N__23326),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__3334 (
            .O(N__23323),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__3333 (
            .O(N__23316),
            .I(N__23311));
    InMux I__3332 (
            .O(N__23315),
            .I(N__23308));
    InMux I__3331 (
            .O(N__23314),
            .I(N__23305));
    LocalMux I__3330 (
            .O(N__23311),
            .I(N__23302));
    LocalMux I__3329 (
            .O(N__23308),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__3328 (
            .O(N__23305),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__3327 (
            .O(N__23302),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__3326 (
            .O(N__23295),
            .I(N__23290));
    InMux I__3325 (
            .O(N__23294),
            .I(N__23287));
    InMux I__3324 (
            .O(N__23293),
            .I(N__23284));
    LocalMux I__3323 (
            .O(N__23290),
            .I(N__23281));
    LocalMux I__3322 (
            .O(N__23287),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__3321 (
            .O(N__23284),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__3320 (
            .O(N__23281),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__3319 (
            .O(N__23274),
            .I(N__23270));
    InMux I__3318 (
            .O(N__23273),
            .I(N__23266));
    LocalMux I__3317 (
            .O(N__23270),
            .I(N__23263));
    InMux I__3316 (
            .O(N__23269),
            .I(N__23260));
    LocalMux I__3315 (
            .O(N__23266),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv12 I__3314 (
            .O(N__23263),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__3313 (
            .O(N__23260),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__3312 (
            .O(N__23253),
            .I(N__23249));
    InMux I__3311 (
            .O(N__23252),
            .I(N__23246));
    LocalMux I__3310 (
            .O(N__23249),
            .I(N__23240));
    LocalMux I__3309 (
            .O(N__23246),
            .I(N__23240));
    InMux I__3308 (
            .O(N__23245),
            .I(N__23237));
    Odrv4 I__3307 (
            .O(N__23240),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__3306 (
            .O(N__23237),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    CascadeMux I__3305 (
            .O(N__23232),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__3304 (
            .O(N__23229),
            .I(N__23225));
    InMux I__3303 (
            .O(N__23228),
            .I(N__23222));
    LocalMux I__3302 (
            .O(N__23225),
            .I(N__23216));
    LocalMux I__3301 (
            .O(N__23222),
            .I(N__23216));
    InMux I__3300 (
            .O(N__23221),
            .I(N__23213));
    Odrv4 I__3299 (
            .O(N__23216),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__3298 (
            .O(N__23213),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__3297 (
            .O(N__23208),
            .I(N__23205));
    LocalMux I__3296 (
            .O(N__23205),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__3295 (
            .O(N__23202),
            .I(N__23198));
    InMux I__3294 (
            .O(N__23201),
            .I(N__23194));
    LocalMux I__3293 (
            .O(N__23198),
            .I(N__23191));
    InMux I__3292 (
            .O(N__23197),
            .I(N__23188));
    LocalMux I__3291 (
            .O(N__23194),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv12 I__3290 (
            .O(N__23191),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__3289 (
            .O(N__23188),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    CascadeMux I__3288 (
            .O(N__23181),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__3287 (
            .O(N__23178),
            .I(N__23175));
    LocalMux I__3286 (
            .O(N__23175),
            .I(N__23170));
    InMux I__3285 (
            .O(N__23174),
            .I(N__23167));
    InMux I__3284 (
            .O(N__23173),
            .I(N__23164));
    Odrv4 I__3283 (
            .O(N__23170),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__3282 (
            .O(N__23167),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__3281 (
            .O(N__23164),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__3280 (
            .O(N__23157),
            .I(N__23145));
    InMux I__3279 (
            .O(N__23156),
            .I(N__23142));
    InMux I__3278 (
            .O(N__23155),
            .I(N__23133));
    InMux I__3277 (
            .O(N__23154),
            .I(N__23133));
    InMux I__3276 (
            .O(N__23153),
            .I(N__23133));
    InMux I__3275 (
            .O(N__23152),
            .I(N__23133));
    InMux I__3274 (
            .O(N__23151),
            .I(N__23124));
    InMux I__3273 (
            .O(N__23150),
            .I(N__23124));
    InMux I__3272 (
            .O(N__23149),
            .I(N__23124));
    InMux I__3271 (
            .O(N__23148),
            .I(N__23124));
    LocalMux I__3270 (
            .O(N__23145),
            .I(N__23119));
    LocalMux I__3269 (
            .O(N__23142),
            .I(N__23119));
    LocalMux I__3268 (
            .O(N__23133),
            .I(N__23116));
    LocalMux I__3267 (
            .O(N__23124),
            .I(N__23113));
    Span4Mux_h I__3266 (
            .O(N__23119),
            .I(N__23110));
    Odrv12 I__3265 (
            .O(N__23116),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__3264 (
            .O(N__23113),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__3263 (
            .O(N__23110),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__3262 (
            .O(N__23103),
            .I(N__23100));
    LocalMux I__3261 (
            .O(N__23100),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3260 (
            .O(N__23097),
            .I(N__23092));
    InMux I__3259 (
            .O(N__23096),
            .I(N__23089));
    InMux I__3258 (
            .O(N__23095),
            .I(N__23085));
    LocalMux I__3257 (
            .O(N__23092),
            .I(N__23082));
    LocalMux I__3256 (
            .O(N__23089),
            .I(N__23079));
    InMux I__3255 (
            .O(N__23088),
            .I(N__23076));
    LocalMux I__3254 (
            .O(N__23085),
            .I(N__23073));
    Span4Mux_h I__3253 (
            .O(N__23082),
            .I(N__23068));
    Span4Mux_h I__3252 (
            .O(N__23079),
            .I(N__23068));
    LocalMux I__3251 (
            .O(N__23076),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv12 I__3250 (
            .O(N__23073),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__3249 (
            .O(N__23068),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__3248 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__3247 (
            .O(N__23058),
            .I(N__23055));
    Odrv4 I__3246 (
            .O(N__23055),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3245 (
            .O(N__23052),
            .I(N__23045));
    InMux I__3244 (
            .O(N__23051),
            .I(N__23045));
    InMux I__3243 (
            .O(N__23050),
            .I(N__23042));
    LocalMux I__3242 (
            .O(N__23045),
            .I(N__23038));
    LocalMux I__3241 (
            .O(N__23042),
            .I(N__23035));
    InMux I__3240 (
            .O(N__23041),
            .I(N__23032));
    Span4Mux_h I__3239 (
            .O(N__23038),
            .I(N__23029));
    Odrv4 I__3238 (
            .O(N__23035),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3237 (
            .O(N__23032),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__3236 (
            .O(N__23029),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__3235 (
            .O(N__23022),
            .I(N__23019));
    LocalMux I__3234 (
            .O(N__23019),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__3233 (
            .O(N__23016),
            .I(N__23013));
    LocalMux I__3232 (
            .O(N__23013),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3231 (
            .O(N__23010),
            .I(N__23007));
    LocalMux I__3230 (
            .O(N__23007),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__3229 (
            .O(N__23004),
            .I(N__23000));
    InMux I__3228 (
            .O(N__23003),
            .I(N__22997));
    InMux I__3227 (
            .O(N__23000),
            .I(N__22993));
    LocalMux I__3226 (
            .O(N__22997),
            .I(N__22989));
    InMux I__3225 (
            .O(N__22996),
            .I(N__22986));
    LocalMux I__3224 (
            .O(N__22993),
            .I(N__22983));
    InMux I__3223 (
            .O(N__22992),
            .I(N__22980));
    Sp12to4 I__3222 (
            .O(N__22989),
            .I(N__22975));
    LocalMux I__3221 (
            .O(N__22986),
            .I(N__22975));
    Odrv4 I__3220 (
            .O(N__22983),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__3219 (
            .O(N__22980),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__3218 (
            .O(N__22975),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__3217 (
            .O(N__22968),
            .I(N__22965));
    InMux I__3216 (
            .O(N__22965),
            .I(N__22962));
    LocalMux I__3215 (
            .O(N__22962),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    CascadeMux I__3214 (
            .O(N__22959),
            .I(N__22953));
    InMux I__3213 (
            .O(N__22958),
            .I(N__22950));
    CascadeMux I__3212 (
            .O(N__22957),
            .I(N__22947));
    CascadeMux I__3211 (
            .O(N__22956),
            .I(N__22944));
    InMux I__3210 (
            .O(N__22953),
            .I(N__22941));
    LocalMux I__3209 (
            .O(N__22950),
            .I(N__22938));
    InMux I__3208 (
            .O(N__22947),
            .I(N__22935));
    InMux I__3207 (
            .O(N__22944),
            .I(N__22932));
    LocalMux I__3206 (
            .O(N__22941),
            .I(N__22929));
    Span4Mux_h I__3205 (
            .O(N__22938),
            .I(N__22926));
    LocalMux I__3204 (
            .O(N__22935),
            .I(N__22923));
    LocalMux I__3203 (
            .O(N__22932),
            .I(N__22918));
    Sp12to4 I__3202 (
            .O(N__22929),
            .I(N__22918));
    Odrv4 I__3201 (
            .O(N__22926),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__3200 (
            .O(N__22923),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv12 I__3199 (
            .O(N__22918),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__3198 (
            .O(N__22911),
            .I(N__22908));
    LocalMux I__3197 (
            .O(N__22908),
            .I(N__22905));
    Span4Mux_v I__3196 (
            .O(N__22905),
            .I(N__22902));
    Odrv4 I__3195 (
            .O(N__22902),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__3194 (
            .O(N__22899),
            .I(N__22896));
    LocalMux I__3193 (
            .O(N__22896),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    CascadeMux I__3192 (
            .O(N__22893),
            .I(N__22890));
    InMux I__3191 (
            .O(N__22890),
            .I(N__22887));
    LocalMux I__3190 (
            .O(N__22887),
            .I(N__22881));
    InMux I__3189 (
            .O(N__22886),
            .I(N__22878));
    InMux I__3188 (
            .O(N__22885),
            .I(N__22875));
    InMux I__3187 (
            .O(N__22884),
            .I(N__22872));
    Odrv4 I__3186 (
            .O(N__22881),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__3185 (
            .O(N__22878),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__3184 (
            .O(N__22875),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__3183 (
            .O(N__22872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__3182 (
            .O(N__22863),
            .I(N__22860));
    InMux I__3181 (
            .O(N__22860),
            .I(N__22857));
    LocalMux I__3180 (
            .O(N__22857),
            .I(N__22854));
    Span4Mux_v I__3179 (
            .O(N__22854),
            .I(N__22848));
    InMux I__3178 (
            .O(N__22853),
            .I(N__22843));
    InMux I__3177 (
            .O(N__22852),
            .I(N__22843));
    InMux I__3176 (
            .O(N__22851),
            .I(N__22840));
    Odrv4 I__3175 (
            .O(N__22848),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__3174 (
            .O(N__22843),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__3173 (
            .O(N__22840),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__3172 (
            .O(N__22833),
            .I(N__22830));
    InMux I__3171 (
            .O(N__22830),
            .I(N__22826));
    CascadeMux I__3170 (
            .O(N__22829),
            .I(N__22823));
    LocalMux I__3169 (
            .O(N__22826),
            .I(N__22818));
    InMux I__3168 (
            .O(N__22823),
            .I(N__22813));
    InMux I__3167 (
            .O(N__22822),
            .I(N__22813));
    InMux I__3166 (
            .O(N__22821),
            .I(N__22810));
    Span4Mux_h I__3165 (
            .O(N__22818),
            .I(N__22805));
    LocalMux I__3164 (
            .O(N__22813),
            .I(N__22805));
    LocalMux I__3163 (
            .O(N__22810),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__3162 (
            .O(N__22805),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__3161 (
            .O(N__22800),
            .I(N__22797));
    InMux I__3160 (
            .O(N__22797),
            .I(N__22794));
    LocalMux I__3159 (
            .O(N__22794),
            .I(N__22791));
    Odrv4 I__3158 (
            .O(N__22791),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3157 (
            .O(N__22788),
            .I(N__22784));
    InMux I__3156 (
            .O(N__22787),
            .I(N__22780));
    LocalMux I__3155 (
            .O(N__22784),
            .I(N__22777));
    InMux I__3154 (
            .O(N__22783),
            .I(N__22774));
    LocalMux I__3153 (
            .O(N__22780),
            .I(N__22770));
    Span4Mux_h I__3152 (
            .O(N__22777),
            .I(N__22765));
    LocalMux I__3151 (
            .O(N__22774),
            .I(N__22765));
    InMux I__3150 (
            .O(N__22773),
            .I(N__22762));
    Span4Mux_h I__3149 (
            .O(N__22770),
            .I(N__22755));
    Span4Mux_h I__3148 (
            .O(N__22765),
            .I(N__22755));
    LocalMux I__3147 (
            .O(N__22762),
            .I(N__22755));
    Odrv4 I__3146 (
            .O(N__22755),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__3145 (
            .O(N__22752),
            .I(N__22749));
    LocalMux I__3144 (
            .O(N__22749),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3143 (
            .O(N__22746),
            .I(N__22743));
    LocalMux I__3142 (
            .O(N__22743),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__3141 (
            .O(N__22740),
            .I(N__22737));
    InMux I__3140 (
            .O(N__22737),
            .I(N__22732));
    InMux I__3139 (
            .O(N__22736),
            .I(N__22729));
    InMux I__3138 (
            .O(N__22735),
            .I(N__22726));
    LocalMux I__3137 (
            .O(N__22732),
            .I(N__22723));
    LocalMux I__3136 (
            .O(N__22729),
            .I(N__22718));
    LocalMux I__3135 (
            .O(N__22726),
            .I(N__22718));
    Span4Mux_s3_h I__3134 (
            .O(N__22723),
            .I(N__22714));
    Span4Mux_h I__3133 (
            .O(N__22718),
            .I(N__22711));
    InMux I__3132 (
            .O(N__22717),
            .I(N__22708));
    Odrv4 I__3131 (
            .O(N__22714),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3130 (
            .O(N__22711),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3129 (
            .O(N__22708),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__3128 (
            .O(N__22701),
            .I(N__22698));
    LocalMux I__3127 (
            .O(N__22698),
            .I(N__22695));
    Odrv4 I__3126 (
            .O(N__22695),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    CascadeMux I__3125 (
            .O(N__22692),
            .I(N__22689));
    InMux I__3124 (
            .O(N__22689),
            .I(N__22685));
    InMux I__3123 (
            .O(N__22688),
            .I(N__22682));
    LocalMux I__3122 (
            .O(N__22685),
            .I(N__22677));
    LocalMux I__3121 (
            .O(N__22682),
            .I(N__22674));
    InMux I__3120 (
            .O(N__22681),
            .I(N__22671));
    InMux I__3119 (
            .O(N__22680),
            .I(N__22668));
    Span4Mux_h I__3118 (
            .O(N__22677),
            .I(N__22665));
    Span4Mux_v I__3117 (
            .O(N__22674),
            .I(N__22658));
    LocalMux I__3116 (
            .O(N__22671),
            .I(N__22658));
    LocalMux I__3115 (
            .O(N__22668),
            .I(N__22658));
    Odrv4 I__3114 (
            .O(N__22665),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__3113 (
            .O(N__22658),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    CascadeMux I__3112 (
            .O(N__22653),
            .I(N__22650));
    InMux I__3111 (
            .O(N__22650),
            .I(N__22647));
    LocalMux I__3110 (
            .O(N__22647),
            .I(N__22644));
    Odrv12 I__3109 (
            .O(N__22644),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__3108 (
            .O(N__22641),
            .I(N__22638));
    InMux I__3107 (
            .O(N__22638),
            .I(N__22635));
    LocalMux I__3106 (
            .O(N__22635),
            .I(N__22632));
    Odrv12 I__3105 (
            .O(N__22632),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__3104 (
            .O(N__22629),
            .I(N__22626));
    LocalMux I__3103 (
            .O(N__22626),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    CascadeMux I__3102 (
            .O(N__22623),
            .I(N__22618));
    InMux I__3101 (
            .O(N__22622),
            .I(N__22615));
    InMux I__3100 (
            .O(N__22621),
            .I(N__22611));
    InMux I__3099 (
            .O(N__22618),
            .I(N__22608));
    LocalMux I__3098 (
            .O(N__22615),
            .I(N__22605));
    InMux I__3097 (
            .O(N__22614),
            .I(N__22602));
    LocalMux I__3096 (
            .O(N__22611),
            .I(N__22599));
    LocalMux I__3095 (
            .O(N__22608),
            .I(N__22596));
    Span4Mux_v I__3094 (
            .O(N__22605),
            .I(N__22591));
    LocalMux I__3093 (
            .O(N__22602),
            .I(N__22591));
    Odrv4 I__3092 (
            .O(N__22599),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__3091 (
            .O(N__22596),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__3090 (
            .O(N__22591),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__3089 (
            .O(N__22584),
            .I(N__22581));
    LocalMux I__3088 (
            .O(N__22581),
            .I(N__22578));
    Span4Mux_v I__3087 (
            .O(N__22578),
            .I(N__22575));
    Odrv4 I__3086 (
            .O(N__22575),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__3085 (
            .O(N__22572),
            .I(N__22567));
    InMux I__3084 (
            .O(N__22571),
            .I(N__22564));
    InMux I__3083 (
            .O(N__22570),
            .I(N__22561));
    InMux I__3082 (
            .O(N__22567),
            .I(N__22558));
    LocalMux I__3081 (
            .O(N__22564),
            .I(N__22554));
    LocalMux I__3080 (
            .O(N__22561),
            .I(N__22551));
    LocalMux I__3079 (
            .O(N__22558),
            .I(N__22548));
    InMux I__3078 (
            .O(N__22557),
            .I(N__22545));
    Span4Mux_v I__3077 (
            .O(N__22554),
            .I(N__22542));
    Span4Mux_h I__3076 (
            .O(N__22551),
            .I(N__22539));
    Span4Mux_v I__3075 (
            .O(N__22548),
            .I(N__22534));
    LocalMux I__3074 (
            .O(N__22545),
            .I(N__22534));
    Odrv4 I__3073 (
            .O(N__22542),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3072 (
            .O(N__22539),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__3071 (
            .O(N__22534),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__3070 (
            .O(N__22527),
            .I(N__22524));
    LocalMux I__3069 (
            .O(N__22524),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3068 (
            .O(N__22521),
            .I(N__22517));
    CascadeMux I__3067 (
            .O(N__22520),
            .I(N__22513));
    LocalMux I__3066 (
            .O(N__22517),
            .I(N__22510));
    InMux I__3065 (
            .O(N__22516),
            .I(N__22506));
    InMux I__3064 (
            .O(N__22513),
            .I(N__22503));
    Span4Mux_v I__3063 (
            .O(N__22510),
            .I(N__22500));
    InMux I__3062 (
            .O(N__22509),
            .I(N__22497));
    LocalMux I__3061 (
            .O(N__22506),
            .I(N__22492));
    LocalMux I__3060 (
            .O(N__22503),
            .I(N__22492));
    Odrv4 I__3059 (
            .O(N__22500),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__3058 (
            .O(N__22497),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__3057 (
            .O(N__22492),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__3056 (
            .O(N__22485),
            .I(N__22482));
    LocalMux I__3055 (
            .O(N__22482),
            .I(N__22477));
    InMux I__3054 (
            .O(N__22481),
            .I(N__22474));
    InMux I__3053 (
            .O(N__22480),
            .I(N__22470));
    Span4Mux_v I__3052 (
            .O(N__22477),
            .I(N__22467));
    LocalMux I__3051 (
            .O(N__22474),
            .I(N__22464));
    InMux I__3050 (
            .O(N__22473),
            .I(N__22461));
    LocalMux I__3049 (
            .O(N__22470),
            .I(N__22458));
    Odrv4 I__3048 (
            .O(N__22467),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__3047 (
            .O(N__22464),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__3046 (
            .O(N__22461),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__3045 (
            .O(N__22458),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__3044 (
            .O(N__22449),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ));
    InMux I__3043 (
            .O(N__22446),
            .I(N__22442));
    InMux I__3042 (
            .O(N__22445),
            .I(N__22439));
    LocalMux I__3041 (
            .O(N__22442),
            .I(N__22432));
    LocalMux I__3040 (
            .O(N__22439),
            .I(N__22432));
    InMux I__3039 (
            .O(N__22438),
            .I(N__22429));
    InMux I__3038 (
            .O(N__22437),
            .I(N__22426));
    Span4Mux_h I__3037 (
            .O(N__22432),
            .I(N__22423));
    LocalMux I__3036 (
            .O(N__22429),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__3035 (
            .O(N__22426),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__3034 (
            .O(N__22423),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__3033 (
            .O(N__22416),
            .I(N__22412));
    InMux I__3032 (
            .O(N__22415),
            .I(N__22409));
    LocalMux I__3031 (
            .O(N__22412),
            .I(N__22404));
    LocalMux I__3030 (
            .O(N__22409),
            .I(N__22401));
    InMux I__3029 (
            .O(N__22408),
            .I(N__22398));
    InMux I__3028 (
            .O(N__22407),
            .I(N__22395));
    Span4Mux_v I__3027 (
            .O(N__22404),
            .I(N__22392));
    Span4Mux_v I__3026 (
            .O(N__22401),
            .I(N__22385));
    LocalMux I__3025 (
            .O(N__22398),
            .I(N__22385));
    LocalMux I__3024 (
            .O(N__22395),
            .I(N__22385));
    Span4Mux_v I__3023 (
            .O(N__22392),
            .I(N__22382));
    Span4Mux_v I__3022 (
            .O(N__22385),
            .I(N__22379));
    Odrv4 I__3021 (
            .O(N__22382),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__3020 (
            .O(N__22379),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__3019 (
            .O(N__22374),
            .I(N__22371));
    InMux I__3018 (
            .O(N__22371),
            .I(N__22367));
    InMux I__3017 (
            .O(N__22370),
            .I(N__22363));
    LocalMux I__3016 (
            .O(N__22367),
            .I(N__22360));
    CascadeMux I__3015 (
            .O(N__22366),
            .I(N__22357));
    LocalMux I__3014 (
            .O(N__22363),
            .I(N__22353));
    Span12Mux_s5_h I__3013 (
            .O(N__22360),
            .I(N__22350));
    InMux I__3012 (
            .O(N__22357),
            .I(N__22347));
    InMux I__3011 (
            .O(N__22356),
            .I(N__22344));
    Span4Mux_v I__3010 (
            .O(N__22353),
            .I(N__22341));
    Odrv12 I__3009 (
            .O(N__22350),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3008 (
            .O(N__22347),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__3007 (
            .O(N__22344),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__3006 (
            .O(N__22341),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CascadeMux I__3005 (
            .O(N__22332),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ));
    InMux I__3004 (
            .O(N__22329),
            .I(N__22326));
    LocalMux I__3003 (
            .O(N__22326),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    InMux I__3002 (
            .O(N__22323),
            .I(N__22320));
    LocalMux I__3001 (
            .O(N__22320),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ));
    InMux I__3000 (
            .O(N__22317),
            .I(N__22314));
    LocalMux I__2999 (
            .O(N__22314),
            .I(N__22311));
    Odrv4 I__2998 (
            .O(N__22311),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__2997 (
            .O(N__22308),
            .I(N__22305));
    LocalMux I__2996 (
            .O(N__22305),
            .I(N__22302));
    Odrv4 I__2995 (
            .O(N__22302),
            .I(\current_shift_inst.PI_CTRL.N_167 ));
    InMux I__2994 (
            .O(N__22299),
            .I(N__22296));
    LocalMux I__2993 (
            .O(N__22296),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    InMux I__2992 (
            .O(N__22293),
            .I(N__22290));
    LocalMux I__2991 (
            .O(N__22290),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__2990 (
            .O(N__22287),
            .I(\current_shift_inst.PI_CTRL.N_171_cascade_ ));
    InMux I__2989 (
            .O(N__22284),
            .I(N__22281));
    LocalMux I__2988 (
            .O(N__22281),
            .I(N__22275));
    InMux I__2987 (
            .O(N__22280),
            .I(N__22270));
    InMux I__2986 (
            .O(N__22279),
            .I(N__22270));
    InMux I__2985 (
            .O(N__22278),
            .I(N__22267));
    Span4Mux_v I__2984 (
            .O(N__22275),
            .I(N__22262));
    LocalMux I__2983 (
            .O(N__22270),
            .I(N__22262));
    LocalMux I__2982 (
            .O(N__22267),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2981 (
            .O(N__22262),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__2980 (
            .O(N__22257),
            .I(N__22254));
    InMux I__2979 (
            .O(N__22254),
            .I(N__22251));
    LocalMux I__2978 (
            .O(N__22251),
            .I(N__22248));
    Span4Mux_h I__2977 (
            .O(N__22248),
            .I(N__22245));
    Odrv4 I__2976 (
            .O(N__22245),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__2975 (
            .O(N__22242),
            .I(N__22239));
    InMux I__2974 (
            .O(N__22239),
            .I(N__22235));
    InMux I__2973 (
            .O(N__22238),
            .I(N__22232));
    LocalMux I__2972 (
            .O(N__22235),
            .I(N__22227));
    LocalMux I__2971 (
            .O(N__22232),
            .I(N__22224));
    InMux I__2970 (
            .O(N__22231),
            .I(N__22221));
    InMux I__2969 (
            .O(N__22230),
            .I(N__22218));
    Span4Mux_v I__2968 (
            .O(N__22227),
            .I(N__22215));
    Span4Mux_v I__2967 (
            .O(N__22224),
            .I(N__22208));
    LocalMux I__2966 (
            .O(N__22221),
            .I(N__22208));
    LocalMux I__2965 (
            .O(N__22218),
            .I(N__22208));
    Odrv4 I__2964 (
            .O(N__22215),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__2963 (
            .O(N__22208),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__2962 (
            .O(N__22203),
            .I(N__22200));
    LocalMux I__2961 (
            .O(N__22200),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__2960 (
            .O(N__22197),
            .I(N__22193));
    InMux I__2959 (
            .O(N__22196),
            .I(N__22189));
    InMux I__2958 (
            .O(N__22193),
            .I(N__22185));
    InMux I__2957 (
            .O(N__22192),
            .I(N__22182));
    LocalMux I__2956 (
            .O(N__22189),
            .I(N__22179));
    CascadeMux I__2955 (
            .O(N__22188),
            .I(N__22176));
    LocalMux I__2954 (
            .O(N__22185),
            .I(N__22173));
    LocalMux I__2953 (
            .O(N__22182),
            .I(N__22168));
    Span4Mux_h I__2952 (
            .O(N__22179),
            .I(N__22168));
    InMux I__2951 (
            .O(N__22176),
            .I(N__22165));
    Odrv4 I__2950 (
            .O(N__22173),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__2949 (
            .O(N__22168),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__2948 (
            .O(N__22165),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__2947 (
            .O(N__22158),
            .I(N__22155));
    LocalMux I__2946 (
            .O(N__22155),
            .I(N__22152));
    Span4Mux_h I__2945 (
            .O(N__22152),
            .I(N__22149));
    Odrv4 I__2944 (
            .O(N__22149),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__2943 (
            .O(N__22146),
            .I(N__22142));
    InMux I__2942 (
            .O(N__22145),
            .I(N__22139));
    InMux I__2941 (
            .O(N__22142),
            .I(N__22135));
    LocalMux I__2940 (
            .O(N__22139),
            .I(N__22131));
    InMux I__2939 (
            .O(N__22138),
            .I(N__22128));
    LocalMux I__2938 (
            .O(N__22135),
            .I(N__22125));
    InMux I__2937 (
            .O(N__22134),
            .I(N__22122));
    Span4Mux_h I__2936 (
            .O(N__22131),
            .I(N__22119));
    LocalMux I__2935 (
            .O(N__22128),
            .I(N__22116));
    Span4Mux_v I__2934 (
            .O(N__22125),
            .I(N__22111));
    LocalMux I__2933 (
            .O(N__22122),
            .I(N__22111));
    Odrv4 I__2932 (
            .O(N__22119),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__2931 (
            .O(N__22116),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__2930 (
            .O(N__22111),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__2929 (
            .O(N__22104),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2928 (
            .O(N__22101),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2927 (
            .O(N__22098),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2926 (
            .O(N__22095),
            .I(bfn_5_7_0_));
    InMux I__2925 (
            .O(N__22092),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2924 (
            .O(N__22089),
            .I(N__22086));
    LocalMux I__2923 (
            .O(N__22086),
            .I(N__22083));
    Span4Mux_v I__2922 (
            .O(N__22083),
            .I(N__22080));
    Odrv4 I__2921 (
            .O(N__22080),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    CascadeMux I__2920 (
            .O(N__22077),
            .I(N__22074));
    InMux I__2919 (
            .O(N__22074),
            .I(N__22071));
    LocalMux I__2918 (
            .O(N__22071),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__2917 (
            .O(N__22068),
            .I(N__22065));
    LocalMux I__2916 (
            .O(N__22065),
            .I(N__22060));
    InMux I__2915 (
            .O(N__22064),
            .I(N__22057));
    InMux I__2914 (
            .O(N__22063),
            .I(N__22053));
    Span12Mux_s4_h I__2913 (
            .O(N__22060),
            .I(N__22048));
    LocalMux I__2912 (
            .O(N__22057),
            .I(N__22048));
    InMux I__2911 (
            .O(N__22056),
            .I(N__22045));
    LocalMux I__2910 (
            .O(N__22053),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__2909 (
            .O(N__22048),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__2908 (
            .O(N__22045),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__2907 (
            .O(N__22038),
            .I(N__22034));
    InMux I__2906 (
            .O(N__22037),
            .I(N__22030));
    InMux I__2905 (
            .O(N__22034),
            .I(N__22027));
    InMux I__2904 (
            .O(N__22033),
            .I(N__22024));
    LocalMux I__2903 (
            .O(N__22030),
            .I(counterZ0Z_1));
    LocalMux I__2902 (
            .O(N__22027),
            .I(counterZ0Z_1));
    LocalMux I__2901 (
            .O(N__22024),
            .I(counterZ0Z_1));
    InMux I__2900 (
            .O(N__22017),
            .I(N__22009));
    InMux I__2899 (
            .O(N__22016),
            .I(N__22009));
    InMux I__2898 (
            .O(N__22015),
            .I(N__22006));
    InMux I__2897 (
            .O(N__22014),
            .I(N__22003));
    LocalMux I__2896 (
            .O(N__22009),
            .I(counterZ0Z_0));
    LocalMux I__2895 (
            .O(N__22006),
            .I(counterZ0Z_0));
    LocalMux I__2894 (
            .O(N__22003),
            .I(counterZ0Z_0));
    InMux I__2893 (
            .O(N__21996),
            .I(N__21989));
    InMux I__2892 (
            .O(N__21995),
            .I(N__21989));
    InMux I__2891 (
            .O(N__21994),
            .I(N__21981));
    LocalMux I__2890 (
            .O(N__21989),
            .I(N__21978));
    InMux I__2889 (
            .O(N__21988),
            .I(N__21973));
    InMux I__2888 (
            .O(N__21987),
            .I(N__21973));
    InMux I__2887 (
            .O(N__21986),
            .I(N__21970));
    InMux I__2886 (
            .O(N__21985),
            .I(N__21965));
    InMux I__2885 (
            .O(N__21984),
            .I(N__21965));
    LocalMux I__2884 (
            .O(N__21981),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0 ));
    Odrv4 I__2883 (
            .O(N__21978),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0 ));
    LocalMux I__2882 (
            .O(N__21973),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0 ));
    LocalMux I__2881 (
            .O(N__21970),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0 ));
    LocalMux I__2880 (
            .O(N__21965),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0 ));
    InMux I__2879 (
            .O(N__21954),
            .I(N__21950));
    InMux I__2878 (
            .O(N__21953),
            .I(N__21947));
    LocalMux I__2877 (
            .O(N__21950),
            .I(clk_10khz_i));
    LocalMux I__2876 (
            .O(N__21947),
            .I(clk_10khz_i));
    InMux I__2875 (
            .O(N__21942),
            .I(bfn_5_6_0_));
    InMux I__2874 (
            .O(N__21939),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2873 (
            .O(N__21936),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2872 (
            .O(N__21933),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2871 (
            .O(N__21930),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2870 (
            .O(N__21927),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    InMux I__2869 (
            .O(N__21924),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    InMux I__2868 (
            .O(N__21921),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    InMux I__2867 (
            .O(N__21918),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__2866 (
            .O(N__21915),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__2865 (
            .O(N__21912),
            .I(N__21908));
    InMux I__2864 (
            .O(N__21911),
            .I(N__21905));
    LocalMux I__2863 (
            .O(N__21908),
            .I(N__21902));
    LocalMux I__2862 (
            .O(N__21905),
            .I(counterZ0Z_11));
    Odrv4 I__2861 (
            .O(N__21902),
            .I(counterZ0Z_11));
    InMux I__2860 (
            .O(N__21897),
            .I(N__21893));
    InMux I__2859 (
            .O(N__21896),
            .I(N__21890));
    LocalMux I__2858 (
            .O(N__21893),
            .I(counterZ0Z_6));
    LocalMux I__2857 (
            .O(N__21890),
            .I(counterZ0Z_6));
    CascadeMux I__2856 (
            .O(N__21885),
            .I(N__21881));
    InMux I__2855 (
            .O(N__21884),
            .I(N__21878));
    InMux I__2854 (
            .O(N__21881),
            .I(N__21875));
    LocalMux I__2853 (
            .O(N__21878),
            .I(counterZ0Z_12));
    LocalMux I__2852 (
            .O(N__21875),
            .I(counterZ0Z_12));
    InMux I__2851 (
            .O(N__21870),
            .I(N__21866));
    InMux I__2850 (
            .O(N__21869),
            .I(N__21863));
    LocalMux I__2849 (
            .O(N__21866),
            .I(counterZ0Z_10));
    LocalMux I__2848 (
            .O(N__21863),
            .I(counterZ0Z_10));
    CascadeMux I__2847 (
            .O(N__21858),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0Z_1_cascade_ ));
    InMux I__2846 (
            .O(N__21855),
            .I(N__21851));
    InMux I__2845 (
            .O(N__21854),
            .I(N__21848));
    LocalMux I__2844 (
            .O(N__21851),
            .I(counterZ0Z_8));
    LocalMux I__2843 (
            .O(N__21848),
            .I(counterZ0Z_8));
    InMux I__2842 (
            .O(N__21843),
            .I(N__21839));
    InMux I__2841 (
            .O(N__21842),
            .I(N__21836));
    LocalMux I__2840 (
            .O(N__21839),
            .I(counterZ0Z_7));
    LocalMux I__2839 (
            .O(N__21836),
            .I(counterZ0Z_7));
    CascadeMux I__2838 (
            .O(N__21831),
            .I(N__21828));
    InMux I__2837 (
            .O(N__21828),
            .I(N__21824));
    InMux I__2836 (
            .O(N__21827),
            .I(N__21821));
    LocalMux I__2835 (
            .O(N__21824),
            .I(N__21818));
    LocalMux I__2834 (
            .O(N__21821),
            .I(counterZ0Z_9));
    Odrv4 I__2833 (
            .O(N__21818),
            .I(counterZ0Z_9));
    InMux I__2832 (
            .O(N__21813),
            .I(N__21809));
    InMux I__2831 (
            .O(N__21812),
            .I(N__21806));
    LocalMux I__2830 (
            .O(N__21809),
            .I(counterZ0Z_5));
    LocalMux I__2829 (
            .O(N__21806),
            .I(counterZ0Z_5));
    InMux I__2828 (
            .O(N__21801),
            .I(N__21798));
    LocalMux I__2827 (
            .O(N__21798),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0Z_8 ));
    InMux I__2826 (
            .O(N__21795),
            .I(N__21791));
    InMux I__2825 (
            .O(N__21794),
            .I(N__21788));
    LocalMux I__2824 (
            .O(N__21791),
            .I(counterZ0Z_2));
    LocalMux I__2823 (
            .O(N__21788),
            .I(counterZ0Z_2));
    InMux I__2822 (
            .O(N__21783),
            .I(N__21779));
    InMux I__2821 (
            .O(N__21782),
            .I(N__21776));
    LocalMux I__2820 (
            .O(N__21779),
            .I(counterZ0Z_3));
    LocalMux I__2819 (
            .O(N__21776),
            .I(counterZ0Z_3));
    CascadeMux I__2818 (
            .O(N__21771),
            .I(N__21767));
    InMux I__2817 (
            .O(N__21770),
            .I(N__21764));
    InMux I__2816 (
            .O(N__21767),
            .I(N__21761));
    LocalMux I__2815 (
            .O(N__21764),
            .I(counterZ0Z_4));
    LocalMux I__2814 (
            .O(N__21761),
            .I(counterZ0Z_4));
    InMux I__2813 (
            .O(N__21756),
            .I(N__21753));
    LocalMux I__2812 (
            .O(N__21753),
            .I(\current_shift_inst.PI_CTRL.un2_counterZ0Z_7 ));
    InMux I__2811 (
            .O(N__21750),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    InMux I__2810 (
            .O(N__21747),
            .I(N__21744));
    LocalMux I__2809 (
            .O(N__21744),
            .I(N__21741));
    Odrv4 I__2808 (
            .O(N__21741),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__2807 (
            .O(N__21738),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__2806 (
            .O(N__21735),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    InMux I__2805 (
            .O(N__21732),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    InMux I__2804 (
            .O(N__21729),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    InMux I__2803 (
            .O(N__21726),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    InMux I__2802 (
            .O(N__21723),
            .I(N__21720));
    LocalMux I__2801 (
            .O(N__21720),
            .I(N__21717));
    Span4Mux_v I__2800 (
            .O(N__21717),
            .I(N__21714));
    Odrv4 I__2799 (
            .O(N__21714),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__2798 (
            .O(N__21711),
            .I(bfn_4_16_0_));
    InMux I__2797 (
            .O(N__21708),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ));
    InMux I__2796 (
            .O(N__21705),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    InMux I__2795 (
            .O(N__21702),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    InMux I__2794 (
            .O(N__21699),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    InMux I__2793 (
            .O(N__21696),
            .I(N__21693));
    LocalMux I__2792 (
            .O(N__21693),
            .I(N__21690));
    Odrv4 I__2791 (
            .O(N__21690),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__2790 (
            .O(N__21687),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    InMux I__2789 (
            .O(N__21684),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__2788 (
            .O(N__21681),
            .I(N__21675));
    InMux I__2787 (
            .O(N__21680),
            .I(N__21675));
    LocalMux I__2786 (
            .O(N__21675),
            .I(N__21671));
    InMux I__2785 (
            .O(N__21674),
            .I(N__21667));
    Span4Mux_h I__2784 (
            .O(N__21671),
            .I(N__21664));
    InMux I__2783 (
            .O(N__21670),
            .I(N__21661));
    LocalMux I__2782 (
            .O(N__21667),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__2781 (
            .O(N__21664),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__2780 (
            .O(N__21661),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__2779 (
            .O(N__21654),
            .I(N__21651));
    LocalMux I__2778 (
            .O(N__21651),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__2777 (
            .O(N__21648),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    InMux I__2776 (
            .O(N__21645),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    InMux I__2775 (
            .O(N__21642),
            .I(bfn_4_15_0_));
    InMux I__2774 (
            .O(N__21639),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ));
    InMux I__2773 (
            .O(N__21636),
            .I(N__21633));
    LocalMux I__2772 (
            .O(N__21633),
            .I(N__21630));
    Odrv12 I__2771 (
            .O(N__21630),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__2770 (
            .O(N__21627),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ));
    InMux I__2769 (
            .O(N__21624),
            .I(N__21621));
    LocalMux I__2768 (
            .O(N__21621),
            .I(N__21618));
    Span4Mux_h I__2767 (
            .O(N__21618),
            .I(N__21613));
    InMux I__2766 (
            .O(N__21617),
            .I(N__21610));
    InMux I__2765 (
            .O(N__21616),
            .I(N__21607));
    Odrv4 I__2764 (
            .O(N__21613),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__2763 (
            .O(N__21610),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__2762 (
            .O(N__21607),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__2761 (
            .O(N__21600),
            .I(N__21597));
    LocalMux I__2760 (
            .O(N__21597),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__2759 (
            .O(N__21594),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    InMux I__2758 (
            .O(N__21591),
            .I(N__21586));
    InMux I__2757 (
            .O(N__21590),
            .I(N__21580));
    InMux I__2756 (
            .O(N__21589),
            .I(N__21580));
    LocalMux I__2755 (
            .O(N__21586),
            .I(N__21577));
    InMux I__2754 (
            .O(N__21585),
            .I(N__21574));
    LocalMux I__2753 (
            .O(N__21580),
            .I(N__21569));
    Span4Mux_h I__2752 (
            .O(N__21577),
            .I(N__21569));
    LocalMux I__2751 (
            .O(N__21574),
            .I(N__21566));
    Odrv4 I__2750 (
            .O(N__21569),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__2749 (
            .O(N__21566),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__2748 (
            .O(N__21561),
            .I(N__21558));
    LocalMux I__2747 (
            .O(N__21558),
            .I(N__21555));
    Odrv12 I__2746 (
            .O(N__21555),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__2745 (
            .O(N__21552),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    InMux I__2744 (
            .O(N__21549),
            .I(N__21546));
    LocalMux I__2743 (
            .O(N__21546),
            .I(N__21543));
    Span4Mux_h I__2742 (
            .O(N__21543),
            .I(N__21537));
    InMux I__2741 (
            .O(N__21542),
            .I(N__21534));
    InMux I__2740 (
            .O(N__21541),
            .I(N__21529));
    InMux I__2739 (
            .O(N__21540),
            .I(N__21529));
    Odrv4 I__2738 (
            .O(N__21537),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__2737 (
            .O(N__21534),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__2736 (
            .O(N__21529),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__2735 (
            .O(N__21522),
            .I(N__21519));
    LocalMux I__2734 (
            .O(N__21519),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__2733 (
            .O(N__21516),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__2732 (
            .O(N__21513),
            .I(N__21510));
    LocalMux I__2731 (
            .O(N__21510),
            .I(N__21507));
    Span4Mux_v I__2730 (
            .O(N__21507),
            .I(N__21501));
    InMux I__2729 (
            .O(N__21506),
            .I(N__21498));
    InMux I__2728 (
            .O(N__21505),
            .I(N__21493));
    InMux I__2727 (
            .O(N__21504),
            .I(N__21493));
    Odrv4 I__2726 (
            .O(N__21501),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__2725 (
            .O(N__21498),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__2724 (
            .O(N__21493),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__2723 (
            .O(N__21486),
            .I(N__21483));
    LocalMux I__2722 (
            .O(N__21483),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__2721 (
            .O(N__21480),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    InMux I__2720 (
            .O(N__21477),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    InMux I__2719 (
            .O(N__21474),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    InMux I__2718 (
            .O(N__21471),
            .I(bfn_4_14_0_));
    CascadeMux I__2717 (
            .O(N__21468),
            .I(N__21464));
    InMux I__2716 (
            .O(N__21467),
            .I(N__21457));
    InMux I__2715 (
            .O(N__21464),
            .I(N__21457));
    InMux I__2714 (
            .O(N__21463),
            .I(N__21454));
    InMux I__2713 (
            .O(N__21462),
            .I(N__21451));
    LocalMux I__2712 (
            .O(N__21457),
            .I(N__21448));
    LocalMux I__2711 (
            .O(N__21454),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__2710 (
            .O(N__21451),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__2709 (
            .O(N__21448),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__2708 (
            .O(N__21441),
            .I(N__21438));
    LocalMux I__2707 (
            .O(N__21438),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__2706 (
            .O(N__21435),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ));
    InMux I__2705 (
            .O(N__21432),
            .I(N__21429));
    LocalMux I__2704 (
            .O(N__21429),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    InMux I__2703 (
            .O(N__21426),
            .I(N__21423));
    LocalMux I__2702 (
            .O(N__21423),
            .I(N__21418));
    InMux I__2701 (
            .O(N__21422),
            .I(N__21414));
    InMux I__2700 (
            .O(N__21421),
            .I(N__21411));
    Span4Mux_v I__2699 (
            .O(N__21418),
            .I(N__21408));
    InMux I__2698 (
            .O(N__21417),
            .I(N__21405));
    LocalMux I__2697 (
            .O(N__21414),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__2696 (
            .O(N__21411),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    Odrv4 I__2695 (
            .O(N__21408),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__2694 (
            .O(N__21405),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    CascadeMux I__2693 (
            .O(N__21396),
            .I(N__21393));
    InMux I__2692 (
            .O(N__21393),
            .I(N__21390));
    LocalMux I__2691 (
            .O(N__21390),
            .I(N__21387));
    Odrv4 I__2690 (
            .O(N__21387),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__2689 (
            .O(N__21384),
            .I(N__21381));
    LocalMux I__2688 (
            .O(N__21381),
            .I(N__21378));
    Span4Mux_v I__2687 (
            .O(N__21378),
            .I(N__21373));
    InMux I__2686 (
            .O(N__21377),
            .I(N__21370));
    InMux I__2685 (
            .O(N__21376),
            .I(N__21367));
    Odrv4 I__2684 (
            .O(N__21373),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2683 (
            .O(N__21370),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2682 (
            .O(N__21367),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__2681 (
            .O(N__21360),
            .I(N__21357));
    LocalMux I__2680 (
            .O(N__21357),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__2679 (
            .O(N__21354),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2678 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__2677 (
            .O(N__21348),
            .I(N__21345));
    Span12Mux_s6_v I__2676 (
            .O(N__21345),
            .I(N__21342));
    Span12Mux_h I__2675 (
            .O(N__21342),
            .I(N__21339));
    Odrv12 I__2674 (
            .O(N__21339),
            .I(pwm_output_c));
    CascadeMux I__2673 (
            .O(N__21336),
            .I(\current_shift_inst.PI_CTRL.N_170_cascade_ ));
    CascadeMux I__2672 (
            .O(N__21333),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    InMux I__2671 (
            .O(N__21330),
            .I(N__21327));
    LocalMux I__2670 (
            .O(N__21327),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    InMux I__2669 (
            .O(N__21324),
            .I(N__21321));
    LocalMux I__2668 (
            .O(N__21321),
            .I(\current_shift_inst.PI_CTRL.N_168 ));
    CascadeMux I__2667 (
            .O(N__21318),
            .I(N__21315));
    InMux I__2666 (
            .O(N__21315),
            .I(N__21312));
    LocalMux I__2665 (
            .O(N__21312),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    InMux I__2664 (
            .O(N__21309),
            .I(N__21306));
    LocalMux I__2663 (
            .O(N__21306),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    CascadeMux I__2662 (
            .O(N__21303),
            .I(N__21300));
    InMux I__2661 (
            .O(N__21300),
            .I(N__21297));
    LocalMux I__2660 (
            .O(N__21297),
            .I(N__21294));
    Odrv4 I__2659 (
            .O(N__21294),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    InMux I__2658 (
            .O(N__21291),
            .I(N__21288));
    LocalMux I__2657 (
            .O(N__21288),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2656 (
            .O(N__21285),
            .I(N__21282));
    InMux I__2655 (
            .O(N__21282),
            .I(N__21279));
    LocalMux I__2654 (
            .O(N__21279),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    InMux I__2653 (
            .O(N__21276),
            .I(N__21273));
    LocalMux I__2652 (
            .O(N__21273),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2651 (
            .O(N__21270),
            .I(N__21267));
    InMux I__2650 (
            .O(N__21267),
            .I(N__21264));
    LocalMux I__2649 (
            .O(N__21264),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    InMux I__2648 (
            .O(N__21261),
            .I(N__21258));
    LocalMux I__2647 (
            .O(N__21258),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2646 (
            .O(N__21255),
            .I(N__21252));
    LocalMux I__2645 (
            .O(N__21252),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    CascadeMux I__2644 (
            .O(N__21249),
            .I(N__21246));
    InMux I__2643 (
            .O(N__21246),
            .I(N__21243));
    LocalMux I__2642 (
            .O(N__21243),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2641 (
            .O(N__21240),
            .I(N__21237));
    InMux I__2640 (
            .O(N__21237),
            .I(N__21234));
    LocalMux I__2639 (
            .O(N__21234),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2638 (
            .O(N__21231),
            .I(N__21228));
    LocalMux I__2637 (
            .O(N__21228),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2636 (
            .O(N__21225),
            .I(N__21222));
    InMux I__2635 (
            .O(N__21222),
            .I(N__21219));
    LocalMux I__2634 (
            .O(N__21219),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    InMux I__2633 (
            .O(N__21216),
            .I(N__21213));
    LocalMux I__2632 (
            .O(N__21213),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2631 (
            .O(N__21210),
            .I(N__21207));
    InMux I__2630 (
            .O(N__21207),
            .I(N__21204));
    LocalMux I__2629 (
            .O(N__21204),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2628 (
            .O(N__21201),
            .I(N__21198));
    LocalMux I__2627 (
            .O(N__21198),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2626 (
            .O(N__21195),
            .I(N__21192));
    InMux I__2625 (
            .O(N__21192),
            .I(N__21189));
    LocalMux I__2624 (
            .O(N__21189),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2623 (
            .O(N__21186),
            .I(N__21183));
    LocalMux I__2622 (
            .O(N__21183),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2621 (
            .O(N__21180),
            .I(un5_counter_cry_6));
    InMux I__2620 (
            .O(N__21177),
            .I(un5_counter_cry_7));
    InMux I__2619 (
            .O(N__21174),
            .I(bfn_3_19_0_));
    InMux I__2618 (
            .O(N__21171),
            .I(un5_counter_cry_9));
    InMux I__2617 (
            .O(N__21168),
            .I(un5_counter_cry_10));
    InMux I__2616 (
            .O(N__21165),
            .I(un5_counter_cry_11));
    CascadeMux I__2615 (
            .O(N__21162),
            .I(N__21159));
    InMux I__2614 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__2613 (
            .O(N__21156),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__2612 (
            .O(N__21153),
            .I(N__21150));
    LocalMux I__2611 (
            .O(N__21150),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2610 (
            .O(N__21147),
            .I(N__21144));
    InMux I__2609 (
            .O(N__21144),
            .I(N__21141));
    LocalMux I__2608 (
            .O(N__21141),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    InMux I__2607 (
            .O(N__21138),
            .I(N__21135));
    LocalMux I__2606 (
            .O(N__21135),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2605 (
            .O(N__21132),
            .I(N__21126));
    CascadeMux I__2604 (
            .O(N__21131),
            .I(N__21122));
    CascadeMux I__2603 (
            .O(N__21130),
            .I(N__21118));
    InMux I__2602 (
            .O(N__21129),
            .I(N__21102));
    InMux I__2601 (
            .O(N__21126),
            .I(N__21102));
    InMux I__2600 (
            .O(N__21125),
            .I(N__21102));
    InMux I__2599 (
            .O(N__21122),
            .I(N__21102));
    InMux I__2598 (
            .O(N__21121),
            .I(N__21102));
    InMux I__2597 (
            .O(N__21118),
            .I(N__21102));
    InMux I__2596 (
            .O(N__21117),
            .I(N__21102));
    LocalMux I__2595 (
            .O(N__21102),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__2594 (
            .O(N__21099),
            .I(N__21096));
    LocalMux I__2593 (
            .O(N__21096),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    CascadeMux I__2592 (
            .O(N__21093),
            .I(N__21090));
    InMux I__2591 (
            .O(N__21090),
            .I(N__21087));
    LocalMux I__2590 (
            .O(N__21087),
            .I(N__21084));
    Odrv4 I__2589 (
            .O(N__21084),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__2588 (
            .O(N__21081),
            .I(un5_counter_cry_1));
    InMux I__2587 (
            .O(N__21078),
            .I(un5_counter_cry_2));
    InMux I__2586 (
            .O(N__21075),
            .I(un5_counter_cry_3));
    InMux I__2585 (
            .O(N__21072),
            .I(un5_counter_cry_4));
    InMux I__2584 (
            .O(N__21069),
            .I(un5_counter_cry_5));
    InMux I__2583 (
            .O(N__21066),
            .I(N__21063));
    LocalMux I__2582 (
            .O(N__21063),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__2581 (
            .O(N__21060),
            .I(N__21057));
    LocalMux I__2580 (
            .O(N__21057),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    CascadeMux I__2579 (
            .O(N__21054),
            .I(N__21051));
    InMux I__2578 (
            .O(N__21051),
            .I(N__21048));
    LocalMux I__2577 (
            .O(N__21048),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    CascadeMux I__2576 (
            .O(N__21045),
            .I(N__21042));
    InMux I__2575 (
            .O(N__21042),
            .I(N__21039));
    LocalMux I__2574 (
            .O(N__21039),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__2573 (
            .O(N__21036),
            .I(N__21033));
    InMux I__2572 (
            .O(N__21033),
            .I(N__21030));
    LocalMux I__2571 (
            .O(N__21030),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    CascadeMux I__2570 (
            .O(N__21027),
            .I(N__21024));
    InMux I__2569 (
            .O(N__21024),
            .I(N__21021));
    LocalMux I__2568 (
            .O(N__21021),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    CascadeMux I__2567 (
            .O(N__21018),
            .I(N__21015));
    InMux I__2566 (
            .O(N__21015),
            .I(N__21012));
    LocalMux I__2565 (
            .O(N__21012),
            .I(N__21009));
    Odrv4 I__2564 (
            .O(N__21009),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__2563 (
            .O(N__21006),
            .I(N__21003));
    LocalMux I__2562 (
            .O(N__21003),
            .I(N__21000));
    Odrv4 I__2561 (
            .O(N__21000),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    CascadeMux I__2560 (
            .O(N__20997),
            .I(N__20994));
    InMux I__2559 (
            .O(N__20994),
            .I(N__20991));
    LocalMux I__2558 (
            .O(N__20991),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    CascadeMux I__2557 (
            .O(N__20988),
            .I(N__20985));
    InMux I__2556 (
            .O(N__20985),
            .I(N__20982));
    LocalMux I__2555 (
            .O(N__20982),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2554 (
            .O(N__20979),
            .I(N__20976));
    LocalMux I__2553 (
            .O(N__20976),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__2552 (
            .O(N__20973),
            .I(N__20970));
    InMux I__2551 (
            .O(N__20970),
            .I(N__20967));
    LocalMux I__2550 (
            .O(N__20967),
            .I(N__20964));
    Odrv4 I__2549 (
            .O(N__20964),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__2548 (
            .O(N__20961),
            .I(N__20958));
    InMux I__2547 (
            .O(N__20958),
            .I(N__20955));
    LocalMux I__2546 (
            .O(N__20955),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2545 (
            .O(N__20952),
            .I(N__20949));
    LocalMux I__2544 (
            .O(N__20949),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__2543 (
            .O(N__20946),
            .I(N__20943));
    InMux I__2542 (
            .O(N__20943),
            .I(N__20940));
    LocalMux I__2541 (
            .O(N__20940),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__2540 (
            .O(N__20937),
            .I(N__20934));
    InMux I__2539 (
            .O(N__20934),
            .I(N__20931));
    LocalMux I__2538 (
            .O(N__20931),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__2537 (
            .O(N__20928),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    CascadeMux I__2536 (
            .O(N__20925),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__2535 (
            .O(N__20922),
            .I(N__20919));
    InMux I__2534 (
            .O(N__20919),
            .I(N__20916));
    LocalMux I__2533 (
            .O(N__20916),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    InMux I__2532 (
            .O(N__20913),
            .I(N__20910));
    LocalMux I__2531 (
            .O(N__20910),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    CascadeMux I__2530 (
            .O(N__20907),
            .I(N__20904));
    InMux I__2529 (
            .O(N__20904),
            .I(N__20901));
    LocalMux I__2528 (
            .O(N__20901),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__2527 (
            .O(N__20898),
            .I(N__20895));
    InMux I__2526 (
            .O(N__20895),
            .I(N__20892));
    LocalMux I__2525 (
            .O(N__20892),
            .I(N__20889));
    Odrv4 I__2524 (
            .O(N__20889),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2523 (
            .O(N__20886),
            .I(N__20883));
    InMux I__2522 (
            .O(N__20883),
            .I(N__20880));
    LocalMux I__2521 (
            .O(N__20880),
            .I(N__20877));
    Odrv4 I__2520 (
            .O(N__20877),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2519 (
            .O(N__20874),
            .I(N__20870));
    InMux I__2518 (
            .O(N__20873),
            .I(N__20866));
    LocalMux I__2517 (
            .O(N__20870),
            .I(N__20863));
    InMux I__2516 (
            .O(N__20869),
            .I(N__20860));
    LocalMux I__2515 (
            .O(N__20866),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    Odrv12 I__2514 (
            .O(N__20863),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2513 (
            .O(N__20860),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    CascadeMux I__2512 (
            .O(N__20853),
            .I(N__20850));
    InMux I__2511 (
            .O(N__20850),
            .I(N__20847));
    LocalMux I__2510 (
            .O(N__20847),
            .I(N__20844));
    Odrv4 I__2509 (
            .O(N__20844),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__2508 (
            .O(N__20841),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    CascadeMux I__2507 (
            .O(N__20838),
            .I(N__20833));
    InMux I__2506 (
            .O(N__20837),
            .I(N__20830));
    InMux I__2505 (
            .O(N__20836),
            .I(N__20827));
    InMux I__2504 (
            .O(N__20833),
            .I(N__20824));
    LocalMux I__2503 (
            .O(N__20830),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2502 (
            .O(N__20827),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2501 (
            .O(N__20824),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__2500 (
            .O(N__20817),
            .I(N__20814));
    LocalMux I__2499 (
            .O(N__20814),
            .I(N__20811));
    Span4Mux_s3_h I__2498 (
            .O(N__20811),
            .I(N__20808));
    Odrv4 I__2497 (
            .O(N__20808),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__2496 (
            .O(N__20805),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__2495 (
            .O(N__20802),
            .I(N__20797));
    InMux I__2494 (
            .O(N__20801),
            .I(N__20794));
    InMux I__2493 (
            .O(N__20800),
            .I(N__20791));
    LocalMux I__2492 (
            .O(N__20797),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__2491 (
            .O(N__20794),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    LocalMux I__2490 (
            .O(N__20791),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    CascadeMux I__2489 (
            .O(N__20784),
            .I(N__20781));
    InMux I__2488 (
            .O(N__20781),
            .I(N__20778));
    LocalMux I__2487 (
            .O(N__20778),
            .I(N__20775));
    Odrv4 I__2486 (
            .O(N__20775),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__2485 (
            .O(N__20772),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__2484 (
            .O(N__20769),
            .I(N__20765));
    InMux I__2483 (
            .O(N__20768),
            .I(N__20762));
    LocalMux I__2482 (
            .O(N__20765),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__2481 (
            .O(N__20762),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__2480 (
            .O(N__20757),
            .I(N__20754));
    LocalMux I__2479 (
            .O(N__20754),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__2478 (
            .O(N__20751),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__2477 (
            .O(N__20748),
            .I(N__20743));
    InMux I__2476 (
            .O(N__20747),
            .I(N__20740));
    InMux I__2475 (
            .O(N__20746),
            .I(N__20737));
    LocalMux I__2474 (
            .O(N__20743),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2473 (
            .O(N__20740),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2472 (
            .O(N__20737),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__2471 (
            .O(N__20730),
            .I(N__20727));
    LocalMux I__2470 (
            .O(N__20727),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__2469 (
            .O(N__20724),
            .I(bfn_3_11_0_));
    InMux I__2468 (
            .O(N__20721),
            .I(N__20717));
    InMux I__2467 (
            .O(N__20720),
            .I(N__20714));
    LocalMux I__2466 (
            .O(N__20717),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2465 (
            .O(N__20714),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__2464 (
            .O(N__20709),
            .I(N__20706));
    LocalMux I__2463 (
            .O(N__20706),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__2462 (
            .O(N__20703),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__2461 (
            .O(N__20700),
            .I(N__20696));
    InMux I__2460 (
            .O(N__20699),
            .I(N__20693));
    LocalMux I__2459 (
            .O(N__20696),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__2458 (
            .O(N__20693),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2457 (
            .O(N__20688),
            .I(N__20685));
    LocalMux I__2456 (
            .O(N__20685),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__2455 (
            .O(N__20682),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__2454 (
            .O(N__20679),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__2453 (
            .O(N__20676),
            .I(N__20673));
    LocalMux I__2452 (
            .O(N__20673),
            .I(N__20670));
    Span4Mux_s3_h I__2451 (
            .O(N__20670),
            .I(N__20667));
    Odrv4 I__2450 (
            .O(N__20667),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__2449 (
            .O(N__20664),
            .I(N__20661));
    LocalMux I__2448 (
            .O(N__20661),
            .I(N__20658));
    Span4Mux_h I__2447 (
            .O(N__20658),
            .I(N__20655));
    Odrv4 I__2446 (
            .O(N__20655),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__2445 (
            .O(N__20652),
            .I(N__20649));
    LocalMux I__2444 (
            .O(N__20649),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__2443 (
            .O(N__20646),
            .I(N__20643));
    LocalMux I__2442 (
            .O(N__20643),
            .I(N__20640));
    Span4Mux_h I__2441 (
            .O(N__20640),
            .I(N__20637));
    Odrv4 I__2440 (
            .O(N__20637),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__2439 (
            .O(N__20634),
            .I(N__20631));
    LocalMux I__2438 (
            .O(N__20631),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__2437 (
            .O(N__20628),
            .I(N__20625));
    LocalMux I__2436 (
            .O(N__20625),
            .I(N__20622));
    Span4Mux_h I__2435 (
            .O(N__20622),
            .I(N__20619));
    Odrv4 I__2434 (
            .O(N__20619),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2433 (
            .O(N__20616),
            .I(N__20613));
    LocalMux I__2432 (
            .O(N__20613),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__2431 (
            .O(N__20610),
            .I(N__20607));
    LocalMux I__2430 (
            .O(N__20607),
            .I(N__20604));
    Span4Mux_v I__2429 (
            .O(N__20604),
            .I(N__20601));
    Odrv4 I__2428 (
            .O(N__20601),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2427 (
            .O(N__20598),
            .I(N__20595));
    LocalMux I__2426 (
            .O(N__20595),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__2425 (
            .O(N__20592),
            .I(N__20589));
    LocalMux I__2424 (
            .O(N__20589),
            .I(N__20586));
    Span4Mux_v I__2423 (
            .O(N__20586),
            .I(N__20583));
    Odrv4 I__2422 (
            .O(N__20583),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__2421 (
            .O(N__20580),
            .I(N__20577));
    LocalMux I__2420 (
            .O(N__20577),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__2419 (
            .O(N__20574),
            .I(N__20569));
    InMux I__2418 (
            .O(N__20573),
            .I(N__20566));
    InMux I__2417 (
            .O(N__20572),
            .I(N__20563));
    LocalMux I__2416 (
            .O(N__20569),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__2415 (
            .O(N__20566),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__2414 (
            .O(N__20563),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    CascadeMux I__2413 (
            .O(N__20556),
            .I(N__20553));
    InMux I__2412 (
            .O(N__20553),
            .I(N__20550));
    LocalMux I__2411 (
            .O(N__20550),
            .I(N__20547));
    Odrv4 I__2410 (
            .O(N__20547),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__2409 (
            .O(N__20544),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    CascadeMux I__2408 (
            .O(N__20541),
            .I(N__20537));
    InMux I__2407 (
            .O(N__20540),
            .I(N__20530));
    InMux I__2406 (
            .O(N__20537),
            .I(N__20527));
    InMux I__2405 (
            .O(N__20536),
            .I(N__20522));
    InMux I__2404 (
            .O(N__20535),
            .I(N__20522));
    InMux I__2403 (
            .O(N__20534),
            .I(N__20519));
    InMux I__2402 (
            .O(N__20533),
            .I(N__20510));
    LocalMux I__2401 (
            .O(N__20530),
            .I(N__20503));
    LocalMux I__2400 (
            .O(N__20527),
            .I(N__20503));
    LocalMux I__2399 (
            .O(N__20522),
            .I(N__20503));
    LocalMux I__2398 (
            .O(N__20519),
            .I(N__20500));
    InMux I__2397 (
            .O(N__20518),
            .I(N__20487));
    InMux I__2396 (
            .O(N__20517),
            .I(N__20487));
    InMux I__2395 (
            .O(N__20516),
            .I(N__20487));
    InMux I__2394 (
            .O(N__20515),
            .I(N__20487));
    InMux I__2393 (
            .O(N__20514),
            .I(N__20487));
    InMux I__2392 (
            .O(N__20513),
            .I(N__20487));
    LocalMux I__2391 (
            .O(N__20510),
            .I(N__20480));
    Span4Mux_v I__2390 (
            .O(N__20503),
            .I(N__20480));
    Span4Mux_h I__2389 (
            .O(N__20500),
            .I(N__20480));
    LocalMux I__2388 (
            .O(N__20487),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2387 (
            .O(N__20480),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2386 (
            .O(N__20475),
            .I(N__20472));
    LocalMux I__2385 (
            .O(N__20472),
            .I(N__20468));
    InMux I__2384 (
            .O(N__20471),
            .I(N__20465));
    Span4Mux_h I__2383 (
            .O(N__20468),
            .I(N__20460));
    LocalMux I__2382 (
            .O(N__20465),
            .I(N__20460));
    Odrv4 I__2381 (
            .O(N__20460),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__2380 (
            .O(N__20457),
            .I(N__20454));
    LocalMux I__2379 (
            .O(N__20454),
            .I(N__20451));
    Odrv4 I__2378 (
            .O(N__20451),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2377 (
            .O(N__20448),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    InMux I__2376 (
            .O(N__20445),
            .I(N__20442));
    LocalMux I__2375 (
            .O(N__20442),
            .I(N__20439));
    Odrv12 I__2374 (
            .O(N__20439),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2373 (
            .O(N__20436),
            .I(N__20433));
    LocalMux I__2372 (
            .O(N__20433),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2371 (
            .O(N__20430),
            .I(N__20427));
    LocalMux I__2370 (
            .O(N__20427),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    CascadeMux I__2369 (
            .O(N__20424),
            .I(N__20418));
    CascadeMux I__2368 (
            .O(N__20423),
            .I(N__20415));
    InMux I__2367 (
            .O(N__20422),
            .I(N__20411));
    CascadeMux I__2366 (
            .O(N__20421),
            .I(N__20403));
    InMux I__2365 (
            .O(N__20418),
            .I(N__20398));
    InMux I__2364 (
            .O(N__20415),
            .I(N__20398));
    CascadeMux I__2363 (
            .O(N__20414),
            .I(N__20395));
    LocalMux I__2362 (
            .O(N__20411),
            .I(N__20392));
    InMux I__2361 (
            .O(N__20410),
            .I(N__20389));
    InMux I__2360 (
            .O(N__20409),
            .I(N__20378));
    InMux I__2359 (
            .O(N__20408),
            .I(N__20378));
    InMux I__2358 (
            .O(N__20407),
            .I(N__20378));
    InMux I__2357 (
            .O(N__20406),
            .I(N__20378));
    InMux I__2356 (
            .O(N__20403),
            .I(N__20378));
    LocalMux I__2355 (
            .O(N__20398),
            .I(N__20375));
    InMux I__2354 (
            .O(N__20395),
            .I(N__20372));
    Span4Mux_h I__2353 (
            .O(N__20392),
            .I(N__20369));
    LocalMux I__2352 (
            .O(N__20389),
            .I(N__20366));
    LocalMux I__2351 (
            .O(N__20378),
            .I(N__20363));
    Span4Mux_h I__2350 (
            .O(N__20375),
            .I(N__20358));
    LocalMux I__2349 (
            .O(N__20372),
            .I(N__20358));
    Span4Mux_v I__2348 (
            .O(N__20369),
            .I(N__20355));
    Span4Mux_h I__2347 (
            .O(N__20366),
            .I(N__20352));
    Span4Mux_v I__2346 (
            .O(N__20363),
            .I(N__20347));
    Span4Mux_s2_h I__2345 (
            .O(N__20358),
            .I(N__20347));
    Odrv4 I__2344 (
            .O(N__20355),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2343 (
            .O(N__20352),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2342 (
            .O(N__20347),
            .I(\pwm_generator_inst.N_17 ));
    CascadeMux I__2341 (
            .O(N__20340),
            .I(N__20331));
    InMux I__2340 (
            .O(N__20339),
            .I(N__20324));
    InMux I__2339 (
            .O(N__20338),
            .I(N__20324));
    InMux I__2338 (
            .O(N__20337),
            .I(N__20321));
    InMux I__2337 (
            .O(N__20336),
            .I(N__20318));
    InMux I__2336 (
            .O(N__20335),
            .I(N__20307));
    InMux I__2335 (
            .O(N__20334),
            .I(N__20307));
    InMux I__2334 (
            .O(N__20331),
            .I(N__20307));
    InMux I__2333 (
            .O(N__20330),
            .I(N__20307));
    InMux I__2332 (
            .O(N__20329),
            .I(N__20307));
    LocalMux I__2331 (
            .O(N__20324),
            .I(N__20301));
    LocalMux I__2330 (
            .O(N__20321),
            .I(N__20301));
    LocalMux I__2329 (
            .O(N__20318),
            .I(N__20296));
    LocalMux I__2328 (
            .O(N__20307),
            .I(N__20296));
    InMux I__2327 (
            .O(N__20306),
            .I(N__20293));
    Span4Mux_v I__2326 (
            .O(N__20301),
            .I(N__20290));
    Span4Mux_h I__2325 (
            .O(N__20296),
            .I(N__20285));
    LocalMux I__2324 (
            .O(N__20293),
            .I(N__20285));
    Odrv4 I__2323 (
            .O(N__20290),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2322 (
            .O(N__20285),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2321 (
            .O(N__20280),
            .I(N__20271));
    InMux I__2320 (
            .O(N__20279),
            .I(N__20264));
    InMux I__2319 (
            .O(N__20278),
            .I(N__20264));
    CascadeMux I__2318 (
            .O(N__20277),
            .I(N__20258));
    CascadeMux I__2317 (
            .O(N__20276),
            .I(N__20255));
    CascadeMux I__2316 (
            .O(N__20275),
            .I(N__20252));
    CascadeMux I__2315 (
            .O(N__20274),
            .I(N__20247));
    InMux I__2314 (
            .O(N__20271),
            .I(N__20244));
    InMux I__2313 (
            .O(N__20270),
            .I(N__20239));
    InMux I__2312 (
            .O(N__20269),
            .I(N__20239));
    LocalMux I__2311 (
            .O(N__20264),
            .I(N__20229));
    InMux I__2310 (
            .O(N__20263),
            .I(N__20222));
    InMux I__2309 (
            .O(N__20262),
            .I(N__20222));
    InMux I__2308 (
            .O(N__20261),
            .I(N__20222));
    InMux I__2307 (
            .O(N__20258),
            .I(N__20215));
    InMux I__2306 (
            .O(N__20255),
            .I(N__20215));
    InMux I__2305 (
            .O(N__20252),
            .I(N__20215));
    InMux I__2304 (
            .O(N__20251),
            .I(N__20210));
    InMux I__2303 (
            .O(N__20250),
            .I(N__20210));
    InMux I__2302 (
            .O(N__20247),
            .I(N__20207));
    LocalMux I__2301 (
            .O(N__20244),
            .I(N__20202));
    LocalMux I__2300 (
            .O(N__20239),
            .I(N__20202));
    InMux I__2299 (
            .O(N__20238),
            .I(N__20176));
    InMux I__2298 (
            .O(N__20237),
            .I(N__20176));
    InMux I__2297 (
            .O(N__20236),
            .I(N__20176));
    InMux I__2296 (
            .O(N__20235),
            .I(N__20176));
    InMux I__2295 (
            .O(N__20234),
            .I(N__20176));
    InMux I__2294 (
            .O(N__20233),
            .I(N__20176));
    InMux I__2293 (
            .O(N__20232),
            .I(N__20176));
    Span4Mux_s1_h I__2292 (
            .O(N__20229),
            .I(N__20171));
    LocalMux I__2291 (
            .O(N__20222),
            .I(N__20171));
    LocalMux I__2290 (
            .O(N__20215),
            .I(N__20162));
    LocalMux I__2289 (
            .O(N__20210),
            .I(N__20162));
    LocalMux I__2288 (
            .O(N__20207),
            .I(N__20162));
    Span4Mux_v I__2287 (
            .O(N__20202),
            .I(N__20162));
    InMux I__2286 (
            .O(N__20201),
            .I(N__20157));
    InMux I__2285 (
            .O(N__20200),
            .I(N__20157));
    InMux I__2284 (
            .O(N__20199),
            .I(N__20154));
    InMux I__2283 (
            .O(N__20198),
            .I(N__20137));
    InMux I__2282 (
            .O(N__20197),
            .I(N__20137));
    InMux I__2281 (
            .O(N__20196),
            .I(N__20137));
    InMux I__2280 (
            .O(N__20195),
            .I(N__20137));
    InMux I__2279 (
            .O(N__20194),
            .I(N__20137));
    InMux I__2278 (
            .O(N__20193),
            .I(N__20137));
    InMux I__2277 (
            .O(N__20192),
            .I(N__20137));
    InMux I__2276 (
            .O(N__20191),
            .I(N__20137));
    LocalMux I__2275 (
            .O(N__20176),
            .I(N__20132));
    Span4Mux_v I__2274 (
            .O(N__20171),
            .I(N__20132));
    Odrv4 I__2273 (
            .O(N__20162),
            .I(N_19_1));
    LocalMux I__2272 (
            .O(N__20157),
            .I(N_19_1));
    LocalMux I__2271 (
            .O(N__20154),
            .I(N_19_1));
    LocalMux I__2270 (
            .O(N__20137),
            .I(N_19_1));
    Odrv4 I__2269 (
            .O(N__20132),
            .I(N_19_1));
    InMux I__2268 (
            .O(N__20121),
            .I(N__20118));
    LocalMux I__2267 (
            .O(N__20118),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2266 (
            .O(N__20115),
            .I(N__20112));
    LocalMux I__2265 (
            .O(N__20112),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2264 (
            .O(N__20109),
            .I(N__20106));
    LocalMux I__2263 (
            .O(N__20106),
            .I(N__20103));
    Span4Mux_v I__2262 (
            .O(N__20103),
            .I(N__20100));
    Odrv4 I__2261 (
            .O(N__20100),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__2260 (
            .O(N__20097),
            .I(N__20094));
    LocalMux I__2259 (
            .O(N__20094),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__2258 (
            .O(N__20091),
            .I(N__20088));
    LocalMux I__2257 (
            .O(N__20088),
            .I(N__20085));
    Span4Mux_v I__2256 (
            .O(N__20085),
            .I(N__20082));
    Odrv4 I__2255 (
            .O(N__20082),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__2254 (
            .O(N__20079),
            .I(N__20076));
    LocalMux I__2253 (
            .O(N__20076),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__2252 (
            .O(N__20073),
            .I(N__20070));
    LocalMux I__2251 (
            .O(N__20070),
            .I(N__20067));
    Span4Mux_v I__2250 (
            .O(N__20067),
            .I(N__20064));
    Odrv4 I__2249 (
            .O(N__20064),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__2248 (
            .O(N__20061),
            .I(N__20058));
    LocalMux I__2247 (
            .O(N__20058),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__2246 (
            .O(N__20055),
            .I(N__20052));
    LocalMux I__2245 (
            .O(N__20052),
            .I(N__20049));
    Span4Mux_h I__2244 (
            .O(N__20049),
            .I(N__20046));
    Odrv4 I__2243 (
            .O(N__20046),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__2242 (
            .O(N__20043),
            .I(N__20040));
    LocalMux I__2241 (
            .O(N__20040),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__2240 (
            .O(N__20037),
            .I(N__20034));
    LocalMux I__2239 (
            .O(N__20034),
            .I(N__20031));
    Span4Mux_h I__2238 (
            .O(N__20031),
            .I(N__20028));
    Odrv4 I__2237 (
            .O(N__20028),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__2236 (
            .O(N__20025),
            .I(N__20022));
    LocalMux I__2235 (
            .O(N__20022),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__2234 (
            .O(N__20019),
            .I(N__20016));
    LocalMux I__2233 (
            .O(N__20016),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__2232 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__2231 (
            .O(N__20010),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    InMux I__2230 (
            .O(N__20007),
            .I(N__20004));
    LocalMux I__2229 (
            .O(N__20004),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__2228 (
            .O(N__20001),
            .I(N__19998));
    LocalMux I__2227 (
            .O(N__19998),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2226 (
            .O(N__19995),
            .I(N__19992));
    LocalMux I__2225 (
            .O(N__19992),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__2224 (
            .O(N__19989),
            .I(N__19986));
    LocalMux I__2223 (
            .O(N__19986),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2222 (
            .O(N__19983),
            .I(N__19980));
    LocalMux I__2221 (
            .O(N__19980),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2220 (
            .O(N__19977),
            .I(N__19974));
    LocalMux I__2219 (
            .O(N__19974),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2218 (
            .O(N__19971),
            .I(N__19967));
    InMux I__2217 (
            .O(N__19970),
            .I(N__19964));
    LocalMux I__2216 (
            .O(N__19967),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    LocalMux I__2215 (
            .O(N__19964),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    CascadeMux I__2214 (
            .O(N__19959),
            .I(N__19955));
    InMux I__2213 (
            .O(N__19958),
            .I(N__19952));
    InMux I__2212 (
            .O(N__19955),
            .I(N__19949));
    LocalMux I__2211 (
            .O(N__19952),
            .I(N__19946));
    LocalMux I__2210 (
            .O(N__19949),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    Odrv4 I__2209 (
            .O(N__19946),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    CascadeMux I__2208 (
            .O(N__19941),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__2207 (
            .O(N__19938),
            .I(N__19935));
    LocalMux I__2206 (
            .O(N__19935),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2205 (
            .O(N__19932),
            .I(N__19928));
    InMux I__2204 (
            .O(N__19931),
            .I(N__19925));
    LocalMux I__2203 (
            .O(N__19928),
            .I(N__19920));
    LocalMux I__2202 (
            .O(N__19925),
            .I(N__19920));
    Span4Mux_s3_h I__2201 (
            .O(N__19920),
            .I(N__19917));
    Odrv4 I__2200 (
            .O(N__19917),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2199 (
            .O(N__19914),
            .I(N__19910));
    InMux I__2198 (
            .O(N__19913),
            .I(N__19907));
    LocalMux I__2197 (
            .O(N__19910),
            .I(N__19902));
    LocalMux I__2196 (
            .O(N__19907),
            .I(N__19902));
    Odrv4 I__2195 (
            .O(N__19902),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    CascadeMux I__2194 (
            .O(N__19899),
            .I(N__19896));
    InMux I__2193 (
            .O(N__19896),
            .I(N__19893));
    LocalMux I__2192 (
            .O(N__19893),
            .I(N__19889));
    InMux I__2191 (
            .O(N__19892),
            .I(N__19886));
    Odrv4 I__2190 (
            .O(N__19889),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2189 (
            .O(N__19886),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2188 (
            .O(N__19881),
            .I(N__19878));
    LocalMux I__2187 (
            .O(N__19878),
            .I(N__19874));
    InMux I__2186 (
            .O(N__19877),
            .I(N__19871));
    Odrv4 I__2185 (
            .O(N__19874),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__2184 (
            .O(N__19871),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2183 (
            .O(N__19866),
            .I(N__19863));
    LocalMux I__2182 (
            .O(N__19863),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2181 (
            .O(N__19860),
            .I(N__19857));
    LocalMux I__2180 (
            .O(N__19857),
            .I(N__19854));
    Span12Mux_s11_v I__2179 (
            .O(N__19854),
            .I(N__19851));
    Odrv12 I__2178 (
            .O(N__19851),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2177 (
            .O(N__19848),
            .I(N__19844));
    InMux I__2176 (
            .O(N__19847),
            .I(N__19841));
    LocalMux I__2175 (
            .O(N__19844),
            .I(N__19838));
    LocalMux I__2174 (
            .O(N__19841),
            .I(N__19835));
    Odrv4 I__2173 (
            .O(N__19838),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    Odrv4 I__2172 (
            .O(N__19835),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    CascadeMux I__2171 (
            .O(N__19830),
            .I(N__19827));
    InMux I__2170 (
            .O(N__19827),
            .I(N__19823));
    InMux I__2169 (
            .O(N__19826),
            .I(N__19820));
    LocalMux I__2168 (
            .O(N__19823),
            .I(N__19815));
    LocalMux I__2167 (
            .O(N__19820),
            .I(N__19815));
    Odrv4 I__2166 (
            .O(N__19815),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2165 (
            .O(N__19812),
            .I(N__19808));
    InMux I__2164 (
            .O(N__19811),
            .I(N__19805));
    LocalMux I__2163 (
            .O(N__19808),
            .I(N__19802));
    LocalMux I__2162 (
            .O(N__19805),
            .I(N__19799));
    Span4Mux_v I__2161 (
            .O(N__19802),
            .I(N__19796));
    Odrv4 I__2160 (
            .O(N__19799),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    Odrv4 I__2159 (
            .O(N__19796),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2158 (
            .O(N__19791),
            .I(N__19788));
    LocalMux I__2157 (
            .O(N__19788),
            .I(N__19785));
    Span12Mux_v I__2156 (
            .O(N__19785),
            .I(N__19782));
    Odrv12 I__2155 (
            .O(N__19782),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2154 (
            .O(N__19779),
            .I(N__19775));
    InMux I__2153 (
            .O(N__19778),
            .I(N__19772));
    LocalMux I__2152 (
            .O(N__19775),
            .I(N__19769));
    LocalMux I__2151 (
            .O(N__19772),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    Odrv4 I__2150 (
            .O(N__19769),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2149 (
            .O(N__19764),
            .I(N__19760));
    InMux I__2148 (
            .O(N__19763),
            .I(N__19757));
    LocalMux I__2147 (
            .O(N__19760),
            .I(N__19754));
    LocalMux I__2146 (
            .O(N__19757),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    Odrv4 I__2145 (
            .O(N__19754),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2144 (
            .O(N__19749),
            .I(N__19743));
    InMux I__2143 (
            .O(N__19748),
            .I(N__19743));
    LocalMux I__2142 (
            .O(N__19743),
            .I(N__19740));
    Odrv12 I__2141 (
            .O(N__19740),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2140 (
            .O(N__19737),
            .I(N__19733));
    InMux I__2139 (
            .O(N__19736),
            .I(N__19730));
    LocalMux I__2138 (
            .O(N__19733),
            .I(N__19725));
    LocalMux I__2137 (
            .O(N__19730),
            .I(N__19725));
    Odrv4 I__2136 (
            .O(N__19725),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    CascadeMux I__2135 (
            .O(N__19722),
            .I(N__19718));
    CascadeMux I__2134 (
            .O(N__19721),
            .I(N__19715));
    InMux I__2133 (
            .O(N__19718),
            .I(N__19712));
    InMux I__2132 (
            .O(N__19715),
            .I(N__19709));
    LocalMux I__2131 (
            .O(N__19712),
            .I(N__19704));
    LocalMux I__2130 (
            .O(N__19709),
            .I(N__19704));
    Odrv4 I__2129 (
            .O(N__19704),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2128 (
            .O(N__19701),
            .I(N__19697));
    InMux I__2127 (
            .O(N__19700),
            .I(N__19694));
    LocalMux I__2126 (
            .O(N__19697),
            .I(N__19691));
    LocalMux I__2125 (
            .O(N__19694),
            .I(N__19688));
    Odrv4 I__2124 (
            .O(N__19691),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    Odrv4 I__2123 (
            .O(N__19688),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2122 (
            .O(N__19683),
            .I(N__19679));
    InMux I__2121 (
            .O(N__19682),
            .I(N__19676));
    LocalMux I__2120 (
            .O(N__19679),
            .I(N__19673));
    LocalMux I__2119 (
            .O(N__19676),
            .I(N__19670));
    Odrv4 I__2118 (
            .O(N__19673),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    Odrv12 I__2117 (
            .O(N__19670),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2116 (
            .O(N__19665),
            .I(N__19661));
    InMux I__2115 (
            .O(N__19664),
            .I(N__19658));
    LocalMux I__2114 (
            .O(N__19661),
            .I(N__19655));
    LocalMux I__2113 (
            .O(N__19658),
            .I(N__19652));
    Span4Mux_v I__2112 (
            .O(N__19655),
            .I(N__19649));
    Odrv4 I__2111 (
            .O(N__19652),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    Odrv4 I__2110 (
            .O(N__19649),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    CascadeMux I__2109 (
            .O(N__19644),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2108 (
            .O(N__19641),
            .I(N__19638));
    LocalMux I__2107 (
            .O(N__19638),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2106 (
            .O(N__19635),
            .I(N__19632));
    LocalMux I__2105 (
            .O(N__19632),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    InMux I__2104 (
            .O(N__19629),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2103 (
            .O(N__19626),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2102 (
            .O(N__19623),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2101 (
            .O(N__19620),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2100 (
            .O(N__19617),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2099 (
            .O(N__19614),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2098 (
            .O(N__19611),
            .I(N__19607));
    CascadeMux I__2097 (
            .O(N__19610),
            .I(N__19601));
    LocalMux I__2096 (
            .O(N__19607),
            .I(N__19597));
    InMux I__2095 (
            .O(N__19606),
            .I(N__19594));
    InMux I__2094 (
            .O(N__19605),
            .I(N__19587));
    InMux I__2093 (
            .O(N__19604),
            .I(N__19587));
    InMux I__2092 (
            .O(N__19601),
            .I(N__19587));
    CascadeMux I__2091 (
            .O(N__19600),
            .I(N__19583));
    Span4Mux_v I__2090 (
            .O(N__19597),
            .I(N__19573));
    LocalMux I__2089 (
            .O(N__19594),
            .I(N__19573));
    LocalMux I__2088 (
            .O(N__19587),
            .I(N__19573));
    InMux I__2087 (
            .O(N__19586),
            .I(N__19570));
    InMux I__2086 (
            .O(N__19583),
            .I(N__19561));
    InMux I__2085 (
            .O(N__19582),
            .I(N__19561));
    InMux I__2084 (
            .O(N__19581),
            .I(N__19561));
    InMux I__2083 (
            .O(N__19580),
            .I(N__19561));
    Span4Mux_v I__2082 (
            .O(N__19573),
            .I(N__19558));
    LocalMux I__2081 (
            .O(N__19570),
            .I(N__19553));
    LocalMux I__2080 (
            .O(N__19561),
            .I(N__19553));
    Sp12to4 I__2079 (
            .O(N__19558),
            .I(N__19548));
    Span12Mux_s10_v I__2078 (
            .O(N__19553),
            .I(N__19548));
    Odrv12 I__2077 (
            .O(N__19548),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2076 (
            .O(N__19545),
            .I(N__19542));
    LocalMux I__2075 (
            .O(N__19542),
            .I(N__19538));
    InMux I__2074 (
            .O(N__19541),
            .I(N__19535));
    Odrv4 I__2073 (
            .O(N__19538),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2072 (
            .O(N__19535),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    CascadeMux I__2071 (
            .O(N__19530),
            .I(N__19527));
    InMux I__2070 (
            .O(N__19527),
            .I(N__19523));
    CascadeMux I__2069 (
            .O(N__19526),
            .I(N__19520));
    LocalMux I__2068 (
            .O(N__19523),
            .I(N__19517));
    InMux I__2067 (
            .O(N__19520),
            .I(N__19514));
    Span4Mux_v I__2066 (
            .O(N__19517),
            .I(N__19509));
    LocalMux I__2065 (
            .O(N__19514),
            .I(N__19509));
    Odrv4 I__2064 (
            .O(N__19509),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    CascadeMux I__2063 (
            .O(N__19506),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ));
    InMux I__2062 (
            .O(N__19503),
            .I(N__19498));
    CascadeMux I__2061 (
            .O(N__19502),
            .I(N__19495));
    CascadeMux I__2060 (
            .O(N__19501),
            .I(N__19492));
    LocalMux I__2059 (
            .O(N__19498),
            .I(N__19488));
    InMux I__2058 (
            .O(N__19495),
            .I(N__19481));
    InMux I__2057 (
            .O(N__19492),
            .I(N__19481));
    InMux I__2056 (
            .O(N__19491),
            .I(N__19481));
    Span4Mux_s2_h I__2055 (
            .O(N__19488),
            .I(N__19472));
    LocalMux I__2054 (
            .O(N__19481),
            .I(N__19472));
    InMux I__2053 (
            .O(N__19480),
            .I(N__19469));
    InMux I__2052 (
            .O(N__19479),
            .I(N__19462));
    InMux I__2051 (
            .O(N__19478),
            .I(N__19462));
    InMux I__2050 (
            .O(N__19477),
            .I(N__19462));
    Span4Mux_v I__2049 (
            .O(N__19472),
            .I(N__19459));
    LocalMux I__2048 (
            .O(N__19469),
            .I(N__19454));
    LocalMux I__2047 (
            .O(N__19462),
            .I(N__19454));
    Odrv4 I__2046 (
            .O(N__19459),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv12 I__2045 (
            .O(N__19454),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2044 (
            .O(N__19449),
            .I(N__19446));
    LocalMux I__2043 (
            .O(N__19446),
            .I(N__19442));
    InMux I__2042 (
            .O(N__19445),
            .I(N__19439));
    Span4Mux_v I__2041 (
            .O(N__19442),
            .I(N__19434));
    LocalMux I__2040 (
            .O(N__19439),
            .I(N__19434));
    Odrv4 I__2039 (
            .O(N__19434),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2038 (
            .O(N__19431),
            .I(N__19428));
    LocalMux I__2037 (
            .O(N__19428),
            .I(N__19424));
    InMux I__2036 (
            .O(N__19427),
            .I(N__19421));
    Odrv12 I__2035 (
            .O(N__19424),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2034 (
            .O(N__19421),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2033 (
            .O(N__19416),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2032 (
            .O(N__19413),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2031 (
            .O(N__19410),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2030 (
            .O(N__19407),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2029 (
            .O(N__19404),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2028 (
            .O(N__19401),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2027 (
            .O(N__19398),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2026 (
            .O(N__19395),
            .I(bfn_2_16_0_));
    InMux I__2025 (
            .O(N__19392),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2024 (
            .O(N__19389),
            .I(N__19385));
    InMux I__2023 (
            .O(N__19388),
            .I(N__19382));
    LocalMux I__2022 (
            .O(N__19385),
            .I(N__19378));
    LocalMux I__2021 (
            .O(N__19382),
            .I(N__19375));
    InMux I__2020 (
            .O(N__19381),
            .I(N__19372));
    Span4Mux_v I__2019 (
            .O(N__19378),
            .I(N__19369));
    Span4Mux_v I__2018 (
            .O(N__19375),
            .I(N__19364));
    LocalMux I__2017 (
            .O(N__19372),
            .I(N__19364));
    Odrv4 I__2016 (
            .O(N__19369),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2015 (
            .O(N__19364),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2014 (
            .O(N__19359),
            .I(bfn_2_14_0_));
    InMux I__2013 (
            .O(N__19356),
            .I(N__19351));
    InMux I__2012 (
            .O(N__19355),
            .I(N__19348));
    InMux I__2011 (
            .O(N__19354),
            .I(N__19345));
    LocalMux I__2010 (
            .O(N__19351),
            .I(N__19342));
    LocalMux I__2009 (
            .O(N__19348),
            .I(N__19339));
    LocalMux I__2008 (
            .O(N__19345),
            .I(N__19336));
    Span4Mux_v I__2007 (
            .O(N__19342),
            .I(N__19331));
    Span4Mux_s2_h I__2006 (
            .O(N__19339),
            .I(N__19331));
    Odrv12 I__2005 (
            .O(N__19336),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2004 (
            .O(N__19331),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2003 (
            .O(N__19326),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2002 (
            .O(N__19323),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2001 (
            .O(N__19320),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2000 (
            .O(N__19317),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__1999 (
            .O(N__19314),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__1998 (
            .O(N__19311),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__1997 (
            .O(N__19308),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__1996 (
            .O(N__19305),
            .I(bfn_2_15_0_));
    InMux I__1995 (
            .O(N__19302),
            .I(N__19299));
    LocalMux I__1994 (
            .O(N__19299),
            .I(N__19296));
    Span4Mux_v I__1993 (
            .O(N__19296),
            .I(N__19292));
    InMux I__1992 (
            .O(N__19295),
            .I(N__19289));
    Span4Mux_s2_h I__1991 (
            .O(N__19292),
            .I(N__19286));
    LocalMux I__1990 (
            .O(N__19289),
            .I(N__19283));
    Odrv4 I__1989 (
            .O(N__19286),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    Odrv4 I__1988 (
            .O(N__19283),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__1987 (
            .O(N__19278),
            .I(N__19275));
    LocalMux I__1986 (
            .O(N__19275),
            .I(N__19272));
    Span4Mux_v I__1985 (
            .O(N__19272),
            .I(N__19269));
    Odrv4 I__1984 (
            .O(N__19269),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__1983 (
            .O(N__19266),
            .I(N__19263));
    LocalMux I__1982 (
            .O(N__19263),
            .I(N__19260));
    Span4Mux_v I__1981 (
            .O(N__19260),
            .I(N__19257));
    Odrv4 I__1980 (
            .O(N__19257),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__1979 (
            .O(N__19254),
            .I(N__19251));
    LocalMux I__1978 (
            .O(N__19251),
            .I(N__19248));
    Span4Mux_s3_h I__1977 (
            .O(N__19248),
            .I(N__19245));
    Odrv4 I__1976 (
            .O(N__19245),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__1975 (
            .O(N__19242),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__1974 (
            .O(N__19239),
            .I(N__19236));
    LocalMux I__1973 (
            .O(N__19236),
            .I(N__19233));
    Span4Mux_s3_h I__1972 (
            .O(N__19233),
            .I(N__19230));
    Odrv4 I__1971 (
            .O(N__19230),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__1970 (
            .O(N__19227),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__1969 (
            .O(N__19224),
            .I(N__19219));
    InMux I__1968 (
            .O(N__19223),
            .I(N__19216));
    InMux I__1967 (
            .O(N__19222),
            .I(N__19213));
    LocalMux I__1966 (
            .O(N__19219),
            .I(N__19210));
    LocalMux I__1965 (
            .O(N__19216),
            .I(N__19205));
    LocalMux I__1964 (
            .O(N__19213),
            .I(N__19205));
    Span4Mux_s3_h I__1963 (
            .O(N__19210),
            .I(N__19200));
    Span4Mux_s3_h I__1962 (
            .O(N__19205),
            .I(N__19200));
    Odrv4 I__1961 (
            .O(N__19200),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__1960 (
            .O(N__19197),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__1959 (
            .O(N__19194),
            .I(N__19188));
    InMux I__1958 (
            .O(N__19193),
            .I(N__19183));
    InMux I__1957 (
            .O(N__19192),
            .I(N__19183));
    InMux I__1956 (
            .O(N__19191),
            .I(N__19180));
    LocalMux I__1955 (
            .O(N__19188),
            .I(N__19177));
    LocalMux I__1954 (
            .O(N__19183),
            .I(N__19172));
    LocalMux I__1953 (
            .O(N__19180),
            .I(N__19172));
    Span4Mux_v I__1952 (
            .O(N__19177),
            .I(N__19167));
    Span4Mux_v I__1951 (
            .O(N__19172),
            .I(N__19167));
    Odrv4 I__1950 (
            .O(N__19167),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__1949 (
            .O(N__19164),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__1948 (
            .O(N__19161),
            .I(N__19158));
    InMux I__1947 (
            .O(N__19158),
            .I(N__19153));
    InMux I__1946 (
            .O(N__19157),
            .I(N__19150));
    InMux I__1945 (
            .O(N__19156),
            .I(N__19147));
    LocalMux I__1944 (
            .O(N__19153),
            .I(N__19144));
    LocalMux I__1943 (
            .O(N__19150),
            .I(N__19141));
    LocalMux I__1942 (
            .O(N__19147),
            .I(N__19138));
    Span4Mux_s2_h I__1941 (
            .O(N__19144),
            .I(N__19133));
    Span4Mux_v I__1940 (
            .O(N__19141),
            .I(N__19133));
    Odrv4 I__1939 (
            .O(N__19138),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__1938 (
            .O(N__19133),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__1937 (
            .O(N__19128),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__1936 (
            .O(N__19125),
            .I(N__19120));
    InMux I__1935 (
            .O(N__19124),
            .I(N__19117));
    InMux I__1934 (
            .O(N__19123),
            .I(N__19114));
    LocalMux I__1933 (
            .O(N__19120),
            .I(N__19111));
    LocalMux I__1932 (
            .O(N__19117),
            .I(N__19106));
    LocalMux I__1931 (
            .O(N__19114),
            .I(N__19106));
    Span4Mux_v I__1930 (
            .O(N__19111),
            .I(N__19101));
    Span4Mux_v I__1929 (
            .O(N__19106),
            .I(N__19101));
    Odrv4 I__1928 (
            .O(N__19101),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__1927 (
            .O(N__19098),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__1926 (
            .O(N__19095),
            .I(N__19090));
    InMux I__1925 (
            .O(N__19094),
            .I(N__19087));
    InMux I__1924 (
            .O(N__19093),
            .I(N__19084));
    LocalMux I__1923 (
            .O(N__19090),
            .I(N__19081));
    LocalMux I__1922 (
            .O(N__19087),
            .I(N__19076));
    LocalMux I__1921 (
            .O(N__19084),
            .I(N__19076));
    Span4Mux_v I__1920 (
            .O(N__19081),
            .I(N__19071));
    Span4Mux_v I__1919 (
            .O(N__19076),
            .I(N__19071));
    Odrv4 I__1918 (
            .O(N__19071),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__1917 (
            .O(N__19068),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    CascadeMux I__1916 (
            .O(N__19065),
            .I(N__19062));
    InMux I__1915 (
            .O(N__19062),
            .I(N__19058));
    InMux I__1914 (
            .O(N__19061),
            .I(N__19055));
    LocalMux I__1913 (
            .O(N__19058),
            .I(N__19050));
    LocalMux I__1912 (
            .O(N__19055),
            .I(N__19050));
    Odrv4 I__1911 (
            .O(N__19050),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    InMux I__1910 (
            .O(N__19047),
            .I(N__19044));
    LocalMux I__1909 (
            .O(N__19044),
            .I(N__19041));
    Span4Mux_v I__1908 (
            .O(N__19041),
            .I(N__19038));
    Odrv4 I__1907 (
            .O(N__19038),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    InMux I__1906 (
            .O(N__19035),
            .I(N__19029));
    InMux I__1905 (
            .O(N__19034),
            .I(N__19029));
    LocalMux I__1904 (
            .O(N__19029),
            .I(N__19026));
    Odrv4 I__1903 (
            .O(N__19026),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    CascadeMux I__1902 (
            .O(N__19023),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    InMux I__1901 (
            .O(N__19020),
            .I(N__19017));
    LocalMux I__1900 (
            .O(N__19017),
            .I(N__19014));
    Span4Mux_v I__1899 (
            .O(N__19014),
            .I(N__19011));
    Odrv4 I__1898 (
            .O(N__19011),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__1897 (
            .O(N__19008),
            .I(N__19004));
    InMux I__1896 (
            .O(N__19007),
            .I(N__19001));
    LocalMux I__1895 (
            .O(N__19004),
            .I(N__18996));
    LocalMux I__1894 (
            .O(N__19001),
            .I(N__18996));
    Odrv4 I__1893 (
            .O(N__18996),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    CascadeMux I__1892 (
            .O(N__18993),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ));
    CascadeMux I__1891 (
            .O(N__18990),
            .I(N__18987));
    InMux I__1890 (
            .O(N__18987),
            .I(N__18984));
    LocalMux I__1889 (
            .O(N__18984),
            .I(N__18981));
    Span4Mux_h I__1888 (
            .O(N__18981),
            .I(N__18978));
    Odrv4 I__1887 (
            .O(N__18978),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    CascadeMux I__1886 (
            .O(N__18975),
            .I(N__18972));
    InMux I__1885 (
            .O(N__18972),
            .I(N__18968));
    InMux I__1884 (
            .O(N__18971),
            .I(N__18965));
    LocalMux I__1883 (
            .O(N__18968),
            .I(N__18960));
    LocalMux I__1882 (
            .O(N__18965),
            .I(N__18960));
    Odrv4 I__1881 (
            .O(N__18960),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__1880 (
            .O(N__18957),
            .I(N__18954));
    LocalMux I__1879 (
            .O(N__18954),
            .I(N__18951));
    Odrv12 I__1878 (
            .O(N__18951),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__1877 (
            .O(N__18948),
            .I(N__18945));
    LocalMux I__1876 (
            .O(N__18945),
            .I(N__18941));
    InMux I__1875 (
            .O(N__18944),
            .I(N__18938));
    Span4Mux_h I__1874 (
            .O(N__18941),
            .I(N__18935));
    LocalMux I__1873 (
            .O(N__18938),
            .I(N__18932));
    Odrv4 I__1872 (
            .O(N__18935),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__1871 (
            .O(N__18932),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1870 (
            .O(N__18927),
            .I(N__18924));
    LocalMux I__1869 (
            .O(N__18924),
            .I(N__18921));
    Odrv12 I__1868 (
            .O(N__18921),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    CascadeMux I__1867 (
            .O(N__18918),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__1866 (
            .O(N__18915),
            .I(N__18912));
    LocalMux I__1865 (
            .O(N__18912),
            .I(N__18909));
    Span4Mux_v I__1864 (
            .O(N__18909),
            .I(N__18906));
    Odrv4 I__1863 (
            .O(N__18906),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__1862 (
            .O(N__18903),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ));
    InMux I__1861 (
            .O(N__18900),
            .I(N__18897));
    LocalMux I__1860 (
            .O(N__18897),
            .I(N__18894));
    Span4Mux_h I__1859 (
            .O(N__18894),
            .I(N__18891));
    Odrv4 I__1858 (
            .O(N__18891),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__1857 (
            .O(N__18888),
            .I(N__18885));
    InMux I__1856 (
            .O(N__18885),
            .I(N__18877));
    InMux I__1855 (
            .O(N__18884),
            .I(N__18874));
    InMux I__1854 (
            .O(N__18883),
            .I(N__18867));
    InMux I__1853 (
            .O(N__18882),
            .I(N__18867));
    InMux I__1852 (
            .O(N__18881),
            .I(N__18867));
    InMux I__1851 (
            .O(N__18880),
            .I(N__18864));
    LocalMux I__1850 (
            .O(N__18877),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__1849 (
            .O(N__18874),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__1848 (
            .O(N__18867),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    LocalMux I__1847 (
            .O(N__18864),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    CascadeMux I__1846 (
            .O(N__18855),
            .I(\current_shift_inst.PI_CTRL.N_118_cascade_ ));
    CascadeMux I__1845 (
            .O(N__18852),
            .I(N__18848));
    InMux I__1844 (
            .O(N__18851),
            .I(N__18844));
    InMux I__1843 (
            .O(N__18848),
            .I(N__18839));
    InMux I__1842 (
            .O(N__18847),
            .I(N__18839));
    LocalMux I__1841 (
            .O(N__18844),
            .I(N__18836));
    LocalMux I__1840 (
            .O(N__18839),
            .I(N__18831));
    Span4Mux_v I__1839 (
            .O(N__18836),
            .I(N__18831));
    Odrv4 I__1838 (
            .O(N__18831),
            .I(pwm_duty_input_9));
    InMux I__1837 (
            .O(N__18828),
            .I(N__18822));
    InMux I__1836 (
            .O(N__18827),
            .I(N__18822));
    LocalMux I__1835 (
            .O(N__18822),
            .I(N__18819));
    Odrv4 I__1834 (
            .O(N__18819),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    CascadeMux I__1833 (
            .O(N__18816),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ));
    InMux I__1832 (
            .O(N__18813),
            .I(N__18810));
    LocalMux I__1831 (
            .O(N__18810),
            .I(N__18807));
    Odrv12 I__1830 (
            .O(N__18807),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__1829 (
            .O(N__18804),
            .I(N__18800));
    InMux I__1828 (
            .O(N__18803),
            .I(N__18797));
    LocalMux I__1827 (
            .O(N__18800),
            .I(N__18794));
    LocalMux I__1826 (
            .O(N__18797),
            .I(N__18791));
    Span4Mux_v I__1825 (
            .O(N__18794),
            .I(N__18788));
    Span4Mux_h I__1824 (
            .O(N__18791),
            .I(N__18785));
    Odrv4 I__1823 (
            .O(N__18788),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    Odrv4 I__1822 (
            .O(N__18785),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    CascadeMux I__1821 (
            .O(N__18780),
            .I(N__18777));
    InMux I__1820 (
            .O(N__18777),
            .I(N__18774));
    LocalMux I__1819 (
            .O(N__18774),
            .I(N__18771));
    Span4Mux_v I__1818 (
            .O(N__18771),
            .I(N__18768));
    Odrv4 I__1817 (
            .O(N__18768),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__1816 (
            .O(N__18765),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    InMux I__1815 (
            .O(N__18762),
            .I(N__18759));
    LocalMux I__1814 (
            .O(N__18759),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__1813 (
            .O(N__18756),
            .I(N__18753));
    LocalMux I__1812 (
            .O(N__18753),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    InMux I__1811 (
            .O(N__18750),
            .I(N__18747));
    LocalMux I__1810 (
            .O(N__18747),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    CascadeMux I__1809 (
            .O(N__18744),
            .I(\current_shift_inst.PI_CTRL.N_94_cascade_ ));
    InMux I__1808 (
            .O(N__18741),
            .I(N__18736));
    InMux I__1807 (
            .O(N__18740),
            .I(N__18731));
    InMux I__1806 (
            .O(N__18739),
            .I(N__18731));
    LocalMux I__1805 (
            .O(N__18736),
            .I(\current_shift_inst.PI_CTRL.N_120 ));
    LocalMux I__1804 (
            .O(N__18731),
            .I(\current_shift_inst.PI_CTRL.N_120 ));
    InMux I__1803 (
            .O(N__18726),
            .I(N__18723));
    LocalMux I__1802 (
            .O(N__18723),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__1801 (
            .O(N__18720),
            .I(N__18717));
    InMux I__1800 (
            .O(N__18717),
            .I(N__18713));
    InMux I__1799 (
            .O(N__18716),
            .I(N__18710));
    LocalMux I__1798 (
            .O(N__18713),
            .I(N__18705));
    LocalMux I__1797 (
            .O(N__18710),
            .I(N__18705));
    Span4Mux_h I__1796 (
            .O(N__18705),
            .I(N__18702));
    Span4Mux_v I__1795 (
            .O(N__18702),
            .I(N__18699));
    Odrv4 I__1794 (
            .O(N__18699),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__1793 (
            .O(N__18696),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    InMux I__1792 (
            .O(N__18693),
            .I(N__18689));
    InMux I__1791 (
            .O(N__18692),
            .I(N__18686));
    LocalMux I__1790 (
            .O(N__18689),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    LocalMux I__1789 (
            .O(N__18686),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__1788 (
            .O(N__18681),
            .I(N__18677));
    InMux I__1787 (
            .O(N__18680),
            .I(N__18669));
    InMux I__1786 (
            .O(N__18677),
            .I(N__18669));
    InMux I__1785 (
            .O(N__18676),
            .I(N__18669));
    LocalMux I__1784 (
            .O(N__18669),
            .I(N__18666));
    Span12Mux_h I__1783 (
            .O(N__18666),
            .I(N__18663));
    Odrv12 I__1782 (
            .O(N__18663),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__1781 (
            .O(N__18660),
            .I(N__18657));
    LocalMux I__1780 (
            .O(N__18657),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1779 (
            .O(N__18654),
            .I(N__18651));
    LocalMux I__1778 (
            .O(N__18651),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__1777 (
            .O(N__18648),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__1776 (
            .O(N__18645),
            .I(N__18642));
    LocalMux I__1775 (
            .O(N__18642),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__1774 (
            .O(N__18639),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__1773 (
            .O(N__18636),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__1772 (
            .O(N__18633),
            .I(N__18630));
    LocalMux I__1771 (
            .O(N__18630),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__1770 (
            .O(N__18627),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__1769 (
            .O(N__18624),
            .I(N__18621));
    LocalMux I__1768 (
            .O(N__18621),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__1767 (
            .O(N__18618),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__1766 (
            .O(N__18615),
            .I(N__18612));
    LocalMux I__1765 (
            .O(N__18612),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__1764 (
            .O(N__18609),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__1763 (
            .O(N__18606),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__1762 (
            .O(N__18603),
            .I(bfn_2_8_0_));
    InMux I__1761 (
            .O(N__18600),
            .I(N__18597));
    LocalMux I__1760 (
            .O(N__18597),
            .I(un7_start_stop_0_a3));
    InMux I__1759 (
            .O(N__18594),
            .I(N__18591));
    LocalMux I__1758 (
            .O(N__18591),
            .I(N_34_i_i));
    InMux I__1757 (
            .O(N__18588),
            .I(N__18585));
    LocalMux I__1756 (
            .O(N__18585),
            .I(N__18582));
    Glb2LocalMux I__1755 (
            .O(N__18582),
            .I(N__18579));
    GlobalMux I__1754 (
            .O(N__18579),
            .I(clk_12mhz));
    IoInMux I__1753 (
            .O(N__18576),
            .I(N__18573));
    LocalMux I__1752 (
            .O(N__18573),
            .I(N__18570));
    IoSpan4Mux I__1751 (
            .O(N__18570),
            .I(N__18567));
    Span4Mux_s0_v I__1750 (
            .O(N__18567),
            .I(N__18564));
    Span4Mux_h I__1749 (
            .O(N__18564),
            .I(N__18561));
    Odrv4 I__1748 (
            .O(N__18561),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__1747 (
            .O(N__18558),
            .I(N__18555));
    LocalMux I__1746 (
            .O(N__18555),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    InMux I__1745 (
            .O(N__18552),
            .I(N__18549));
    LocalMux I__1744 (
            .O(N__18549),
            .I(N__18546));
    Odrv12 I__1743 (
            .O(N__18546),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__1742 (
            .O(N__18543),
            .I(N__18540));
    LocalMux I__1741 (
            .O(N__18540),
            .I(N__18537));
    Odrv12 I__1740 (
            .O(N__18537),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__1739 (
            .O(N__18534),
            .I(N__18531));
    LocalMux I__1738 (
            .O(N__18531),
            .I(N__18528));
    Odrv12 I__1737 (
            .O(N__18528),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1736 (
            .O(N__18525),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1735 (
            .O(N__18522),
            .I(N__18519));
    LocalMux I__1734 (
            .O(N__18519),
            .I(N__18516));
    Odrv4 I__1733 (
            .O(N__18516),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    InMux I__1732 (
            .O(N__18513),
            .I(N__18510));
    LocalMux I__1731 (
            .O(N__18510),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ));
    CascadeMux I__1730 (
            .O(N__18507),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__1729 (
            .O(N__18504),
            .I(N__18501));
    LocalMux I__1728 (
            .O(N__18501),
            .I(N__18498));
    Odrv12 I__1727 (
            .O(N__18498),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1726 (
            .O(N__18495),
            .I(bfn_1_15_0_));
    InMux I__1725 (
            .O(N__18492),
            .I(N__18489));
    LocalMux I__1724 (
            .O(N__18489),
            .I(N__18486));
    Odrv12 I__1723 (
            .O(N__18486),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1722 (
            .O(N__18483),
            .I(N__18480));
    LocalMux I__1721 (
            .O(N__18480),
            .I(N__18477));
    Odrv12 I__1720 (
            .O(N__18477),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1719 (
            .O(N__18474),
            .I(N__18471));
    LocalMux I__1718 (
            .O(N__18471),
            .I(N__18468));
    Odrv12 I__1717 (
            .O(N__18468),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1716 (
            .O(N__18465),
            .I(N__18462));
    LocalMux I__1715 (
            .O(N__18462),
            .I(N__18459));
    Odrv12 I__1714 (
            .O(N__18459),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1713 (
            .O(N__18456),
            .I(N__18453));
    LocalMux I__1712 (
            .O(N__18453),
            .I(N__18450));
    Odrv12 I__1711 (
            .O(N__18450),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1710 (
            .O(N__18447),
            .I(N__18444));
    LocalMux I__1709 (
            .O(N__18444),
            .I(N__18441));
    Odrv4 I__1708 (
            .O(N__18441),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1707 (
            .O(N__18438),
            .I(N__18435));
    LocalMux I__1706 (
            .O(N__18435),
            .I(N__18432));
    Odrv4 I__1705 (
            .O(N__18432),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1704 (
            .O(N__18429),
            .I(N__18426));
    LocalMux I__1703 (
            .O(N__18426),
            .I(N__18423));
    Odrv12 I__1702 (
            .O(N__18423),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1701 (
            .O(N__18420),
            .I(N__18417));
    LocalMux I__1700 (
            .O(N__18417),
            .I(N__18414));
    Span4Mux_h I__1699 (
            .O(N__18414),
            .I(N__18411));
    Odrv4 I__1698 (
            .O(N__18411),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1697 (
            .O(N__18408),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1696 (
            .O(N__18405),
            .I(N__18402));
    LocalMux I__1695 (
            .O(N__18402),
            .I(N__18399));
    Span4Mux_h I__1694 (
            .O(N__18399),
            .I(N__18396));
    Odrv4 I__1693 (
            .O(N__18396),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1692 (
            .O(N__18393),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1691 (
            .O(N__18390),
            .I(N__18387));
    LocalMux I__1690 (
            .O(N__18387),
            .I(N__18384));
    Odrv4 I__1689 (
            .O(N__18384),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1688 (
            .O(N__18381),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1687 (
            .O(N__18378),
            .I(N__18375));
    LocalMux I__1686 (
            .O(N__18375),
            .I(N__18372));
    Odrv12 I__1685 (
            .O(N__18372),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1684 (
            .O(N__18369),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    CascadeMux I__1683 (
            .O(N__18366),
            .I(N__18363));
    InMux I__1682 (
            .O(N__18363),
            .I(N__18360));
    LocalMux I__1681 (
            .O(N__18360),
            .I(N__18357));
    Odrv12 I__1680 (
            .O(N__18357),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1679 (
            .O(N__18354),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    InMux I__1678 (
            .O(N__18351),
            .I(N__18348));
    LocalMux I__1677 (
            .O(N__18348),
            .I(N__18345));
    Odrv4 I__1676 (
            .O(N__18345),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1675 (
            .O(N__18342),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    InMux I__1674 (
            .O(N__18339),
            .I(N__18336));
    LocalMux I__1673 (
            .O(N__18336),
            .I(N__18333));
    Odrv4 I__1672 (
            .O(N__18333),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1671 (
            .O(N__18330),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    CascadeMux I__1670 (
            .O(N__18327),
            .I(N__18324));
    InMux I__1669 (
            .O(N__18324),
            .I(N__18321));
    LocalMux I__1668 (
            .O(N__18321),
            .I(N__18318));
    Span4Mux_v I__1667 (
            .O(N__18318),
            .I(N__18315));
    Odrv4 I__1666 (
            .O(N__18315),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1665 (
            .O(N__18312),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    InMux I__1664 (
            .O(N__18309),
            .I(N__18306));
    LocalMux I__1663 (
            .O(N__18306),
            .I(N__18303));
    Span4Mux_v I__1662 (
            .O(N__18303),
            .I(N__18300));
    Span4Mux_v I__1661 (
            .O(N__18300),
            .I(N__18297));
    Odrv4 I__1660 (
            .O(N__18297),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1659 (
            .O(N__18294),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    CascadeMux I__1658 (
            .O(N__18291),
            .I(N__18288));
    InMux I__1657 (
            .O(N__18288),
            .I(N__18285));
    LocalMux I__1656 (
            .O(N__18285),
            .I(N__18282));
    Span4Mux_v I__1655 (
            .O(N__18282),
            .I(N__18279));
    Odrv4 I__1654 (
            .O(N__18279),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1653 (
            .O(N__18276),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    InMux I__1652 (
            .O(N__18273),
            .I(N__18270));
    LocalMux I__1651 (
            .O(N__18270),
            .I(N__18267));
    Span4Mux_v I__1650 (
            .O(N__18267),
            .I(N__18264));
    Odrv4 I__1649 (
            .O(N__18264),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1648 (
            .O(N__18261),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    CascadeMux I__1647 (
            .O(N__18258),
            .I(N__18255));
    InMux I__1646 (
            .O(N__18255),
            .I(N__18252));
    LocalMux I__1645 (
            .O(N__18252),
            .I(N__18249));
    Span4Mux_v I__1644 (
            .O(N__18249),
            .I(N__18246));
    Span4Mux_s1_h I__1643 (
            .O(N__18246),
            .I(N__18243));
    Odrv4 I__1642 (
            .O(N__18243),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1641 (
            .O(N__18240),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    InMux I__1640 (
            .O(N__18237),
            .I(N__18234));
    LocalMux I__1639 (
            .O(N__18234),
            .I(N__18231));
    Span4Mux_v I__1638 (
            .O(N__18231),
            .I(N__18228));
    Odrv4 I__1637 (
            .O(N__18228),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1636 (
            .O(N__18225),
            .I(N__18222));
    LocalMux I__1635 (
            .O(N__18222),
            .I(N__18218));
    InMux I__1634 (
            .O(N__18221),
            .I(N__18215));
    Span4Mux_v I__1633 (
            .O(N__18218),
            .I(N__18207));
    LocalMux I__1632 (
            .O(N__18215),
            .I(N__18207));
    CascadeMux I__1631 (
            .O(N__18214),
            .I(N__18204));
    CascadeMux I__1630 (
            .O(N__18213),
            .I(N__18200));
    CascadeMux I__1629 (
            .O(N__18212),
            .I(N__18196));
    Span4Mux_v I__1628 (
            .O(N__18207),
            .I(N__18192));
    InMux I__1627 (
            .O(N__18204),
            .I(N__18179));
    InMux I__1626 (
            .O(N__18203),
            .I(N__18179));
    InMux I__1625 (
            .O(N__18200),
            .I(N__18179));
    InMux I__1624 (
            .O(N__18199),
            .I(N__18179));
    InMux I__1623 (
            .O(N__18196),
            .I(N__18179));
    InMux I__1622 (
            .O(N__18195),
            .I(N__18179));
    Odrv4 I__1621 (
            .O(N__18192),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    LocalMux I__1620 (
            .O(N__18179),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    InMux I__1619 (
            .O(N__18174),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1618 (
            .O(N__18171),
            .I(N__18168));
    LocalMux I__1617 (
            .O(N__18168),
            .I(N__18165));
    Odrv12 I__1616 (
            .O(N__18165),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1615 (
            .O(N__18162),
            .I(bfn_1_13_0_));
    InMux I__1614 (
            .O(N__18159),
            .I(N__18156));
    LocalMux I__1613 (
            .O(N__18156),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    InMux I__1612 (
            .O(N__18153),
            .I(N__18150));
    LocalMux I__1611 (
            .O(N__18150),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    CascadeMux I__1610 (
            .O(N__18147),
            .I(N__18144));
    InMux I__1609 (
            .O(N__18144),
            .I(N__18141));
    LocalMux I__1608 (
            .O(N__18141),
            .I(N__18138));
    Span4Mux_v I__1607 (
            .O(N__18138),
            .I(N__18135));
    Odrv4 I__1606 (
            .O(N__18135),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    InMux I__1605 (
            .O(N__18132),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1604 (
            .O(N__18129),
            .I(N__18126));
    LocalMux I__1603 (
            .O(N__18126),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    CascadeMux I__1602 (
            .O(N__18123),
            .I(N__18120));
    InMux I__1601 (
            .O(N__18120),
            .I(N__18117));
    LocalMux I__1600 (
            .O(N__18117),
            .I(N__18114));
    Span4Mux_v I__1599 (
            .O(N__18114),
            .I(N__18111));
    Span4Mux_s1_h I__1598 (
            .O(N__18111),
            .I(N__18108));
    Odrv4 I__1597 (
            .O(N__18108),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    InMux I__1596 (
            .O(N__18105),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1595 (
            .O(N__18102),
            .I(N__18099));
    LocalMux I__1594 (
            .O(N__18099),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    CascadeMux I__1593 (
            .O(N__18096),
            .I(N__18093));
    InMux I__1592 (
            .O(N__18093),
            .I(N__18090));
    LocalMux I__1591 (
            .O(N__18090),
            .I(N__18087));
    Span4Mux_v I__1590 (
            .O(N__18087),
            .I(N__18084));
    Odrv4 I__1589 (
            .O(N__18084),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    InMux I__1588 (
            .O(N__18081),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1587 (
            .O(N__18078),
            .I(N__18075));
    LocalMux I__1586 (
            .O(N__18075),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    CascadeMux I__1585 (
            .O(N__18072),
            .I(N__18069));
    InMux I__1584 (
            .O(N__18069),
            .I(N__18066));
    LocalMux I__1583 (
            .O(N__18066),
            .I(N__18063));
    Span4Mux_v I__1582 (
            .O(N__18063),
            .I(N__18060));
    Odrv4 I__1581 (
            .O(N__18060),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    InMux I__1580 (
            .O(N__18057),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1579 (
            .O(N__18054),
            .I(N__18051));
    LocalMux I__1578 (
            .O(N__18051),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    CascadeMux I__1577 (
            .O(N__18048),
            .I(N__18045));
    InMux I__1576 (
            .O(N__18045),
            .I(N__18042));
    LocalMux I__1575 (
            .O(N__18042),
            .I(N__18039));
    Span4Mux_v I__1574 (
            .O(N__18039),
            .I(N__18036));
    Odrv4 I__1573 (
            .O(N__18036),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    InMux I__1572 (
            .O(N__18033),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1571 (
            .O(N__18030),
            .I(N__18027));
    LocalMux I__1570 (
            .O(N__18027),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    CascadeMux I__1569 (
            .O(N__18024),
            .I(N__18021));
    InMux I__1568 (
            .O(N__18021),
            .I(N__18018));
    LocalMux I__1567 (
            .O(N__18018),
            .I(N__18015));
    Span4Mux_v I__1566 (
            .O(N__18015),
            .I(N__18012));
    Odrv4 I__1565 (
            .O(N__18012),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    InMux I__1564 (
            .O(N__18009),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1563 (
            .O(N__18006),
            .I(N__18003));
    LocalMux I__1562 (
            .O(N__18003),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    CascadeMux I__1561 (
            .O(N__18000),
            .I(N__17997));
    InMux I__1560 (
            .O(N__17997),
            .I(N__17994));
    LocalMux I__1559 (
            .O(N__17994),
            .I(N__17991));
    Span4Mux_v I__1558 (
            .O(N__17991),
            .I(N__17988));
    Odrv4 I__1557 (
            .O(N__17988),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    InMux I__1556 (
            .O(N__17985),
            .I(bfn_1_12_0_));
    InMux I__1555 (
            .O(N__17982),
            .I(N__17979));
    LocalMux I__1554 (
            .O(N__17979),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    CascadeMux I__1553 (
            .O(N__17976),
            .I(N__17973));
    InMux I__1552 (
            .O(N__17973),
            .I(N__17970));
    LocalMux I__1551 (
            .O(N__17970),
            .I(N__17967));
    Span4Mux_v I__1550 (
            .O(N__17967),
            .I(N__17964));
    Odrv4 I__1549 (
            .O(N__17964),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    InMux I__1548 (
            .O(N__17961),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    CascadeMux I__1547 (
            .O(N__17958),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    CascadeMux I__1546 (
            .O(N__17955),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ));
    InMux I__1545 (
            .O(N__17952),
            .I(N__17947));
    InMux I__1544 (
            .O(N__17951),
            .I(N__17942));
    InMux I__1543 (
            .O(N__17950),
            .I(N__17942));
    LocalMux I__1542 (
            .O(N__17947),
            .I(N__17939));
    LocalMux I__1541 (
            .O(N__17942),
            .I(pwm_duty_input_6));
    Odrv4 I__1540 (
            .O(N__17939),
            .I(pwm_duty_input_6));
    InMux I__1539 (
            .O(N__17934),
            .I(N__17929));
    InMux I__1538 (
            .O(N__17933),
            .I(N__17924));
    InMux I__1537 (
            .O(N__17932),
            .I(N__17924));
    LocalMux I__1536 (
            .O(N__17929),
            .I(N__17921));
    LocalMux I__1535 (
            .O(N__17924),
            .I(pwm_duty_input_7));
    Odrv4 I__1534 (
            .O(N__17921),
            .I(pwm_duty_input_7));
    InMux I__1533 (
            .O(N__17916),
            .I(N__17911));
    InMux I__1532 (
            .O(N__17915),
            .I(N__17906));
    InMux I__1531 (
            .O(N__17914),
            .I(N__17906));
    LocalMux I__1530 (
            .O(N__17911),
            .I(N__17903));
    LocalMux I__1529 (
            .O(N__17906),
            .I(pwm_duty_input_5));
    Odrv4 I__1528 (
            .O(N__17903),
            .I(pwm_duty_input_5));
    InMux I__1527 (
            .O(N__17898),
            .I(N__17895));
    LocalMux I__1526 (
            .O(N__17895),
            .I(N__17890));
    InMux I__1525 (
            .O(N__17894),
            .I(N__17885));
    InMux I__1524 (
            .O(N__17893),
            .I(N__17885));
    Span4Mux_v I__1523 (
            .O(N__17890),
            .I(N__17882));
    LocalMux I__1522 (
            .O(N__17885),
            .I(pwm_duty_input_4));
    Odrv4 I__1521 (
            .O(N__17882),
            .I(pwm_duty_input_4));
    InMux I__1520 (
            .O(N__17877),
            .I(N__17872));
    InMux I__1519 (
            .O(N__17876),
            .I(N__17869));
    InMux I__1518 (
            .O(N__17875),
            .I(N__17866));
    LocalMux I__1517 (
            .O(N__17872),
            .I(N__17863));
    LocalMux I__1516 (
            .O(N__17869),
            .I(pwm_duty_input_8));
    LocalMux I__1515 (
            .O(N__17866),
            .I(pwm_duty_input_8));
    Odrv4 I__1514 (
            .O(N__17863),
            .I(pwm_duty_input_8));
    CascadeMux I__1513 (
            .O(N__17856),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__1512 (
            .O(N__17853),
            .I(N__17848));
    InMux I__1511 (
            .O(N__17852),
            .I(N__17843));
    InMux I__1510 (
            .O(N__17851),
            .I(N__17843));
    LocalMux I__1509 (
            .O(N__17848),
            .I(N__17840));
    LocalMux I__1508 (
            .O(N__17843),
            .I(pwm_duty_input_3));
    Odrv4 I__1507 (
            .O(N__17840),
            .I(pwm_duty_input_3));
    InMux I__1506 (
            .O(N__17835),
            .I(N__17832));
    LocalMux I__1505 (
            .O(N__17832),
            .I(N__17829));
    Span4Mux_v I__1504 (
            .O(N__17829),
            .I(N__17826));
    Odrv4 I__1503 (
            .O(N__17826),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1502 (
            .O(N__17823),
            .I(N__17820));
    InMux I__1501 (
            .O(N__17820),
            .I(N__17817));
    LocalMux I__1500 (
            .O(N__17817),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    InMux I__1499 (
            .O(N__17814),
            .I(N__17811));
    LocalMux I__1498 (
            .O(N__17811),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    CascadeMux I__1497 (
            .O(N__17808),
            .I(N__17805));
    InMux I__1496 (
            .O(N__17805),
            .I(N__17802));
    LocalMux I__1495 (
            .O(N__17802),
            .I(N__17799));
    Span4Mux_v I__1494 (
            .O(N__17799),
            .I(N__17796));
    Odrv4 I__1493 (
            .O(N__17796),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    InMux I__1492 (
            .O(N__17793),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1491 (
            .O(N__17790),
            .I(N__17786));
    InMux I__1490 (
            .O(N__17789),
            .I(N__17783));
    LocalMux I__1489 (
            .O(N__17786),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1488 (
            .O(N__17783),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    CascadeMux I__1487 (
            .O(N__17778),
            .I(N__17775));
    InMux I__1486 (
            .O(N__17775),
            .I(N__17772));
    LocalMux I__1485 (
            .O(N__17772),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(un5_counter_cry_8),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryinitout(bfn_4_15_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_10_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_11_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_14_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_25_0_));
    defparam IN_MUX_bfv_14_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_26_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_14_26_0_));
    defparam IN_MUX_bfv_14_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_27_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_14_27_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_15 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(\current_shift_inst.control_input_1_cry_23 ),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_2_16_0_));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__39831),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_461_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__31110),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_185_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__28527),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_463_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__34290),
            .CLKHFEN(N__34292),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__34291),
            .RGB2PWM(N__18594),
            .RGB1(rgb_g),
            .CURREN(N__34566),
            .RGB2(rgb_b),
            .RGB1PWM(N__18600),
            .RGB0PWM(N__45622),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_5_4  (
            .in0(N__18225),
            .in1(N__17789),
            .in2(_gnd_net_),
            .in3(N__20199),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19611),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46077),
            .ce(N__24873),
            .sr(N__45526));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_1_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_1_7_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_1_7_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_1_7_4  (
            .in0(N__20201),
            .in1(N__20306),
            .in2(N__20414),
            .in3(N__18762),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46075),
            .ce(),
            .sr(N__45534));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_7_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_7_7 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_7_7  (
            .in0(N__17790),
            .in1(N__20200),
            .in2(N__17778),
            .in3(N__18221),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(N__19266),
            .in2(_gnd_net_),
            .in3(N__18741),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46073),
            .ce(N__24867),
            .sr(N__45541));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_9_0  (
            .in0(N__18740),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19239),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__24824),
            .sr(N__45548));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_9_1 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_9_1  (
            .in0(N__18884),
            .in1(N__18726),
            .in2(N__18720),
            .in3(N__19194),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__24824),
            .sr(N__45548));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_9_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_9_4  (
            .in0(N__19224),
            .in1(N__18750),
            .in2(_gnd_net_),
            .in3(N__18693),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__24824),
            .sr(N__45548));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_9_6 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_9_6  (
            .in0(N__19389),
            .in1(N__19503),
            .in2(N__18888),
            .in3(N__19606),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__24824),
            .sr(N__45548));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_9_7  (
            .in0(N__19254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18739),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46071),
            .ce(N__24824),
            .sr(N__45548));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_0 .LUT_INIT=16'b1010111000001110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_0  (
            .in0(N__19156),
            .in1(N__19491),
            .in2(N__19610),
            .in3(N__18883),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46066),
            .ce(N__24866),
            .sr(N__45555));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_1 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_10_1  (
            .in0(N__18882),
            .in1(N__19605),
            .in2(N__19502),
            .in3(N__19095),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46066),
            .ce(N__24866),
            .sr(N__45555));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_1_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_1_10_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__17932),
            .in2(_gnd_net_),
            .in3(N__17914),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_1_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_1_10_3 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_1_10_3  (
            .in0(N__17875),
            .in1(N__18847),
            .in2(N__17958),
            .in3(N__17950),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_1_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_1_10_4 .LUT_INIT=16'b1111001111110001;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_1_10_4  (
            .in0(N__17852),
            .in1(N__17893),
            .in2(N__17955),
            .in3(N__33147),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_5 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_5  (
            .in0(N__18881),
            .in1(N__19604),
            .in2(N__19501),
            .in3(N__19125),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46066),
            .ce(N__24866),
            .sr(N__45555));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_1_10_6  (
            .in0(N__17951),
            .in1(N__17933),
            .in2(N__18852),
            .in3(N__17915),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_10_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_1_10_7  (
            .in0(N__17894),
            .in1(N__17876),
            .in2(N__17856),
            .in3(N__17851),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__17835),
            .in2(N__17823),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__17814),
            .in2(N__17808),
            .in3(N__17793),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__18153),
            .in2(N__18147),
            .in3(N__18132),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__18129),
            .in2(N__18123),
            .in3(N__18105),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__18102),
            .in2(N__18096),
            .in3(N__18081),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__18078),
            .in2(N__18072),
            .in3(N__18057),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__18054),
            .in2(N__18048),
            .in3(N__18033),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__18030),
            .in2(N__18024),
            .in3(N__18009),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__18006),
            .in2(N__18000),
            .in3(N__17985),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__17982),
            .in2(N__17976),
            .in3(N__17961),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__18195),
            .in2(N__18327),
            .in3(N__18312),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__18309),
            .in2(N__18212),
            .in3(N__18294),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__18199),
            .in2(N__18291),
            .in3(N__18276),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__18273),
            .in2(N__18213),
            .in3(N__18261),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__18203),
            .in2(N__18258),
            .in3(N__18240),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__18237),
            .in2(N__18214),
            .in3(N__18174),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_13_0  (
            .in0(N__18171),
            .in1(N__18522),
            .in2(_gnd_net_),
            .in3(N__18162),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKH62_13_LC_1_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKH62_13_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIKH62_13_LC_1_13_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIKH62_13_LC_1_13_4  (
            .in0(N__19877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19700),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIR3F5_14_LC_1_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIR3F5_14_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIR3F5_14_LC_1_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIR3F5_14_LC_1_13_6  (
            .in0(N__19541),
            .in1(N__19892),
            .in2(N__19530),
            .in3(N__18159),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__20471),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__18420),
            .in2(_gnd_net_),
            .in3(N__18408),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__18405),
            .in2(_gnd_net_),
            .in3(N__18393),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__18390),
            .in2(_gnd_net_),
            .in3(N__18381),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__18378),
            .in2(_gnd_net_),
            .in3(N__18369),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__34449),
            .in2(N__18366),
            .in3(N__18354),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__18351),
            .in2(N__34556),
            .in3(N__18342),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__18339),
            .in2(N__34557),
            .in3(N__18330),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__18504),
            .in2(_gnd_net_),
            .in3(N__18495),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__18492),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__18483),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__18474),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__18465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__18456),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__18447),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__18438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__18429),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__18552),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__18543),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__18534),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18525),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_1_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_1_16_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIV2LD_8_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__19355),
            .in2(_gnd_net_),
            .in3(N__19381),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_16_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_1_16_7  (
            .in0(N__19094),
            .in1(N__19124),
            .in2(N__19161),
            .in3(N__18513),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_11_LC_1_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_11_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_11_LC_1_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNID9E4_11_LC_1_17_2  (
            .in0(N__19914),
            .in1(N__19971),
            .in2(N__19959),
            .in3(N__19932),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_1_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_1_17_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQTKD_5_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__19093),
            .in2(_gnd_net_),
            .in3(N__19157),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_17_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_1_17_4  (
            .in0(N__19356),
            .in1(N__19123),
            .in2(N__18507),
            .in3(N__19388),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_start_stop_0_a3_LC_1_29_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_start_stop_0_a3_LC_1_29_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_start_stop_0_a3_LC_1_29_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_start_stop_0_a3_LC_1_29_5  (
            .in0(_gnd_net_),
            .in1(N__29399),
            .in2(_gnd_net_),
            .in3(N__45620),
            .lcout(un7_start_stop_0_a3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.N_34_i_i_LC_1_30_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.N_34_i_i_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.N_34_i_i_LC_1_30_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.N_34_i_i_LC_1_30_1  (
            .in0(N__45621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29403),
            .lcout(N_34_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_1_30_3.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_1_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_1_30_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_1_30_3 (
            .in0(N__18588),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_2_LC_2_6_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_2_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18558),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(),
            .sr(N__45518));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_6_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_6_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_6_1 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_2_6_1  (
            .in0(N__20409),
            .in1(N__20335),
            .in2(N__20277),
            .in3(N__18615),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(),
            .sr(N__45518));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_2_6_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_2_6_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_2_6_2 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_2_6_2  (
            .in0(N__20250),
            .in1(N__20407),
            .in2(N__20340),
            .in3(N__18633),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(),
            .sr(N__45518));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_6_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_6_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_2_6_3  (
            .in0(N__20406),
            .in1(N__20330),
            .in2(N__20275),
            .in3(N__18645),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(),
            .sr(N__45518));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_2_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_2_6_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_2_6_5 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_2_6_5  (
            .in0(N__18654),
            .in1(N__20251),
            .in2(N__20421),
            .in3(N__20329),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(),
            .sr(N__45518));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_2_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_2_6_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_2_6_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_2_6_7  (
            .in0(N__20408),
            .in1(N__20334),
            .in2(N__20276),
            .in3(N__18624),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46076),
            .ce(),
            .sr(N__45518));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__18927),
            .in2(N__20541),
            .in3(N__20540),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__20457),
            .in2(_gnd_net_),
            .in3(N__18648),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__18756),
            .in2(_gnd_net_),
            .in3(N__18639),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_7_3  (
            .in0(_gnd_net_),
            .in1(N__18957),
            .in2(_gnd_net_),
            .in3(N__18636),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__19278),
            .in2(_gnd_net_),
            .in3(N__18627),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__18813),
            .in2(_gnd_net_),
            .in3(N__18618),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__19047),
            .in2(_gnd_net_),
            .in3(N__18609),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__19020),
            .in2(_gnd_net_),
            .in3(N__18606),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_8_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18990),
            .in3(N__18603),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_8_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_8_1 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_8_1  (
            .in0(N__20676),
            .in1(N__20536),
            .in2(N__18780),
            .in3(N__18765),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_7 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_2_8_7  (
            .in0(N__18804),
            .in1(N__20874),
            .in2(N__20853),
            .in3(N__20535),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_9_0 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_9_0  (
            .in0(N__19478),
            .in1(N__19582),
            .in2(N__18681),
            .in3(N__19192),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(\current_shift_inst.PI_CTRL.N_94_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_9_1 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_9_1  (
            .in0(N__19223),
            .in1(N__18660),
            .in2(N__18744),
            .in3(N__18692),
            .lcout(\current_shift_inst.PI_CTRL.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_9_3 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_9_3  (
            .in0(N__19193),
            .in1(N__18680),
            .in2(N__19600),
            .in3(N__19479),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__19191),
            .in2(_gnd_net_),
            .in3(N__19222),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_9_6 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_9_6  (
            .in0(N__18716),
            .in1(N__19581),
            .in2(N__18696),
            .in3(N__18880),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_9_7  (
            .in0(N__19580),
            .in1(N__18676),
            .in2(_gnd_net_),
            .in3(N__19477),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_23_LC_2_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_23_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_23_LC_2_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPN72_23_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__19682),
            .in2(_gnd_net_),
            .in3(N__19665),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_10_LC_2_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_10_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_10_LC_2_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_10_LC_2_10_1  (
            .in0(N__19860),
            .in1(N__19431),
            .in2(N__18918),
            .in3(N__19449),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_2_10_2  (
            .in0(N__18915),
            .in1(N__19791),
            .in2(N__18903),
            .in3(N__18900),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(\current_shift_inst.PI_CTRL.N_118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_2_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_2_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_2_10_3 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_2_10_3  (
            .in0(N__19586),
            .in1(N__19354),
            .in2(N__18855),
            .in3(N__19480),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46063),
            .ce(N__24872),
            .sr(N__45549));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_11_0  (
            .in0(N__20748),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19061),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_11_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_2_11_2  (
            .in0(N__20574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18944),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_11_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__18827),
            .in2(_gnd_net_),
            .in3(N__20769),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_11_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_11_4  (
            .in0(N__18828),
            .in1(N__20757),
            .in2(N__18816),
            .in3(N__20533),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__18971),
            .in2(_gnd_net_),
            .in3(N__20837),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_11_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_11_6  (
            .in0(N__20873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18803),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_11_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_2_11_7  (
            .in0(N__20802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19295),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_0 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_12_0  (
            .in0(N__20730),
            .in1(N__20747),
            .in2(N__19065),
            .in3(N__20516),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__20721),
            .in2(_gnd_net_),
            .in3(N__19034),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_12_2 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_12_2  (
            .in0(N__19035),
            .in1(N__20709),
            .in2(N__19023),
            .in3(N__20517),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_12_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_12_3  (
            .in0(N__19007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20700),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_12_4  (
            .in0(N__19008),
            .in1(N__20518),
            .in2(N__18993),
            .in3(N__20688),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_12_5 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_12_5  (
            .in0(N__20514),
            .in1(N__20817),
            .in2(N__18975),
            .in3(N__20836),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_2_12_6  (
            .in0(N__20573),
            .in1(N__18948),
            .in2(N__20556),
            .in3(N__20513),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_12_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_12_7 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_12_7  (
            .in0(N__20515),
            .in1(N__20801),
            .in2(N__20784),
            .in3(N__19302),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_2_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_2_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__21426),
            .in2(N__21396),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__21384),
            .in2(N__20973),
            .in3(N__19242),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_2_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_2_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__21624),
            .in2(N__24150),
            .in3(N__19227),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__21591),
            .in2(N__20886),
            .in3(N__19197),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_2_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_2_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__21549),
            .in2(N__20907),
            .in3(N__19164),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_2_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__21513),
            .in2(N__20898),
            .in3(N__19128),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_2_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__22284),
            .in2(N__20988),
            .in3(N__19098),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_2_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__20979),
            .in2(N__22740),
            .in3(N__19068),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__46055),
            .ce(N__24862),
            .sr(N__45565));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_2_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_2_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__23050),
            .in2(N__20937),
            .in3(N__19359),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_2_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__21463),
            .in2(N__20946),
            .in3(N__19326),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_2_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_2_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__21006),
            .in2(N__22863),
            .in3(N__19323),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_2_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_2_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__22196),
            .in2(N__22641),
            .in3(N__19320),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_2_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__22485),
            .in2(N__20961),
            .in3(N__19317),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_2_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__22621),
            .in2(N__21045),
            .in3(N__19314),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_2_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_2_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__21674),
            .in2(N__22653),
            .in3(N__19311),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_2_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_2_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__20952),
            .in2(N__23985),
            .in3(N__19308),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__46047),
            .ce(N__24812),
            .sr(N__45569));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_2_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_2_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__22787),
            .in2(N__21093),
            .in3(N__19305),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_2_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_2_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__21066),
            .in2(N__22374),
            .in3(N__19416),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_2_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_2_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_2_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__22416),
            .in2(N__21054),
            .in3(N__19413),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_2_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_2_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_2_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__22438),
            .in2(N__21027),
            .in3(N__19410),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_2_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_2_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_2_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__21060),
            .in2(N__23004),
            .in3(N__19407),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_2_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_2_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_2_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__23097),
            .in2(N__21018),
            .in3(N__19404),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_2_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_2_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__22521),
            .in2(N__21036),
            .in3(N__19401),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_2_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_2_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_2_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__21099),
            .in2(N__22893),
            .in3(N__19398),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__46039),
            .ce(N__24748),
            .sr(N__45572));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_2_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_2_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_2_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__22068),
            .in2(N__20997),
            .in3(N__19395),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_2_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_2_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_2_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__21117),
            .in2(N__22242),
            .in3(N__19392),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_2_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_2_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_2_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__22571),
            .in2(N__21130),
            .in3(N__19629),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_2_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_2_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_2_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__21121),
            .in2(N__22692),
            .in3(N__19626),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_2_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_2_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_2_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__22958),
            .in2(N__21131),
            .in3(N__19623),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_2_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_2_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_2_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__21125),
            .in2(N__22833),
            .in3(N__19620),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_2_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_2_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_2_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__22145),
            .in2(N__21132),
            .in3(N__19617),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_2_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_2_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_2_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_2_16_7  (
            .in0(N__23579),
            .in1(N__21129),
            .in2(_gnd_net_),
            .in3(N__19614),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46028),
            .ce(N__24786),
            .sr(N__45575));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_2_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_2_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQJB4_15_LC_2_17_0  (
            .in0(N__19545),
            .in1(N__19848),
            .in2(N__19526),
            .in3(N__19811),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_17_1  (
            .in0(N__19866),
            .in1(N__19938),
            .in2(N__19506),
            .in3(N__19635),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_2_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_2_17_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQN62_10_LC_2_17_3  (
            .in0(N__19445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19427),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_2_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_2_17_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5IJ5_27_LC_2_17_4  (
            .in0(N__19970),
            .in1(N__19958),
            .in2(N__19941),
            .in3(N__19826),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_2_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_2_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA3B4_11_LC_2_17_6  (
            .in0(N__19931),
            .in1(N__19913),
            .in2(N__19899),
            .in3(N__19881),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIFF4_21_LC_2_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIFF4_21_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIFF4_21_LC_2_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIFF4_21_LC_2_17_7  (
            .in0(N__19736),
            .in1(N__19778),
            .in2(N__19721),
            .in3(N__19763),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1SC4_17_LC_2_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1SC4_17_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1SC4_17_LC_2_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1SC4_17_LC_2_18_0  (
            .in0(N__19749),
            .in1(N__19847),
            .in2(N__19830),
            .in3(N__19812),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_2_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_2_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNITR72_25_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__19779),
            .in2(_gnd_net_),
            .in3(N__19764),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_2_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_2_18_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFBE4_19_LC_2_18_6  (
            .in0(N__19748),
            .in1(N__19737),
            .in2(N__19722),
            .in3(N__19701),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_2_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_2_18_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI5VT8_23_LC_2_18_7  (
            .in0(N__19683),
            .in1(N__19664),
            .in2(N__19644),
            .in3(N__19641),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_6_LC_3_6_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_3_6_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_3_6_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_3_6_0  (
            .in0(_gnd_net_),
            .in1(N__20019),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_5_LC_3_6_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_3_6_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_3_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_3_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20013),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_7_LC_3_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_3_6_3 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_3_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_3_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19995),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_4_LC_3_6_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_3_6_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_3_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_3_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20007),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_6_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_3_6_5 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_3_6_5  (
            .in0(N__20422),
            .in1(N__20336),
            .in2(N__20274),
            .in3(N__20001),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_0_LC_3_6_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_3_6_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_3_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_3_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19989),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_3_LC_3_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_3_6_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_3_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_3_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20430),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46074),
            .ce(),
            .sr(N__45511));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_7_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_7_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_3_7_0 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_3_7_0  (
            .in0(N__20338),
            .in1(N__19983),
            .in2(N__20423),
            .in3(N__20269),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46072),
            .ce(),
            .sr(N__45519));
    defparam \pwm_generator_inst.threshold_1_LC_3_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_3_7_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_3_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_3_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19977),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46072),
            .ce(),
            .sr(N__45519));
    defparam \pwm_generator_inst.threshold_9_LC_3_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_3_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_3_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_3_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20445),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46072),
            .ce(),
            .sr(N__45519));
    defparam \pwm_generator_inst.threshold_8_LC_3_7_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_3_7_5 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_3_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_3_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20115),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46072),
            .ce(),
            .sr(N__45519));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_7_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_3_7_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_3_7_6  (
            .in0(N__20339),
            .in1(N__20270),
            .in2(N__20424),
            .in3(N__20436),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46072),
            .ce(),
            .sr(N__45519));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_8_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_8_4 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_3_8_4  (
            .in0(N__20410),
            .in1(N__20337),
            .in2(N__20280),
            .in3(N__20121),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46067),
            .ce(),
            .sr(N__45527));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__20097),
            .in2(_gnd_net_),
            .in3(N__20109),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(N__20079),
            .in2(_gnd_net_),
            .in3(N__20091),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__20061),
            .in2(_gnd_net_),
            .in3(N__20073),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__20043),
            .in2(_gnd_net_),
            .in3(N__20055),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__20025),
            .in2(_gnd_net_),
            .in3(N__20037),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__20652),
            .in2(_gnd_net_),
            .in3(N__20664),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__20634),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(N__20616),
            .in2(_gnd_net_),
            .in3(N__20628),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__20598),
            .in2(_gnd_net_),
            .in3(N__20610),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__20580),
            .in2(_gnd_net_),
            .in3(N__20592),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__20572),
            .in2(_gnd_net_),
            .in3(N__20544),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_10_3  (
            .in0(N__20534),
            .in1(N__20475),
            .in2(_gnd_net_),
            .in3(N__20448),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(N__20869),
            .in2(_gnd_net_),
            .in3(N__20841),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20838),
            .in3(N__20805),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(N__20800),
            .in2(_gnd_net_),
            .in3(N__20772),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(N__20768),
            .in2(_gnd_net_),
            .in3(N__20751),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__20746),
            .in2(_gnd_net_),
            .in3(N__20724),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__20720),
            .in2(_gnd_net_),
            .in3(N__20703),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__20699),
            .in2(_gnd_net_),
            .in3(N__20682),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_3_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_3_12_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__22735),
            .in2(_gnd_net_),
            .in3(N__21505),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_3_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_3_12_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_3_12_1  (
            .in0(N__22280),
            .in1(N__23052),
            .in2(N__20928),
            .in3(N__21467),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_3_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_3_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_3_12_2  (
            .in0(N__22736),
            .in1(N__22279),
            .in2(N__21468),
            .in3(N__21504),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_12_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_3_12_3  (
            .in0(N__21589),
            .in1(N__23051),
            .in2(N__20925),
            .in3(N__21540),
            .lcout(\current_shift_inst.PI_CTRL.N_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_3_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_3_12_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_3_12_4  (
            .in0(N__21376),
            .in1(N__21616),
            .in2(_gnd_net_),
            .in3(N__21421),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_3_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_3_12_6 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_3_12_6  (
            .in0(N__21541),
            .in1(N__21590),
            .in2(N__20922),
            .in3(N__20913),
            .lcout(\current_shift_inst.PI_CTRL.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_3_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24029),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(N__24822),
            .sr(N__45561));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24008),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(N__24822),
            .sr(N__45561));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_3_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_3_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24050),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(N__24822),
            .sr(N__45561));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24362),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(N__24822),
            .sr(N__45561));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_3_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_3_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_3_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_3_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24338),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(N__24822),
            .sr(N__45561));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_3_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_3_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24095),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46048),
            .ce(N__24822),
            .sr(N__45561));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_3_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_3_14_1  (
            .in0(N__24221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_2 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_2  (
            .in0(N__21654),
            .in1(N__23900),
            .in2(N__23620),
            .in3(N__23758),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_3 .LUT_INIT=16'b1111001100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_3  (
            .in0(N__23760),
            .in1(N__23603),
            .in2(N__23920),
            .in3(N__21441),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_3_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_3_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_3_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_3_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24549),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24290),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_6 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_3_14_6  (
            .in0(N__21747),
            .in1(N__23901),
            .in2(N__23621),
            .in3(N__23759),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_3_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_3_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24314),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46040),
            .ce(N__24770),
            .sr(N__45566));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_3_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_3_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_3_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24497),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(N__24716),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_3_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_3_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_3_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24431),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(N__24716),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24476),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(N__24716),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_3_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24198),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(N__24716),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24383),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(N__24716),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_3_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24452),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46029),
            .ce(N__24716),
            .sr(N__45570));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_3_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24408),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46018),
            .ce(N__24766),
            .sr(N__45573));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_3_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24267),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46018),
            .ce(N__24766),
            .sr(N__45573));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_3_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_3_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_3_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24941),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46018),
            .ce(N__24766),
            .sr(N__45573));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_3_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_3_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_3_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24915),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46018),
            .ce(N__24766),
            .sr(N__45573));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_3_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_3_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_3_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24971),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46018),
            .ce(N__24766),
            .sr(N__45573));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_3_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_3_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_3_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24527),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46010),
            .ce(N__24703),
            .sr(N__45576));
    defparam un5_counter_cry_1_c_LC_3_18_0.C_ON=1'b1;
    defparam un5_counter_cry_1_c_LC_3_18_0.SEQ_MODE=4'b0000;
    defparam un5_counter_cry_1_c_LC_3_18_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_counter_cry_1_c_LC_3_18_0 (
            .in0(_gnd_net_),
            .in1(N__22015),
            .in2(N__22038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(un5_counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_3_18_1.C_ON=1'b1;
    defparam counter_2_LC_3_18_1.SEQ_MODE=4'b1010;
    defparam counter_2_LC_3_18_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_2_LC_3_18_1 (
            .in0(_gnd_net_),
            .in1(N__21795),
            .in2(_gnd_net_),
            .in3(N__21081),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(un5_counter_cry_1),
            .carryout(un5_counter_cry_2),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_3_LC_3_18_2.C_ON=1'b1;
    defparam counter_3_LC_3_18_2.SEQ_MODE=4'b1010;
    defparam counter_3_LC_3_18_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_3_LC_3_18_2 (
            .in0(_gnd_net_),
            .in1(N__21783),
            .in2(_gnd_net_),
            .in3(N__21078),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(un5_counter_cry_2),
            .carryout(un5_counter_cry_3),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_4_LC_3_18_3.C_ON=1'b1;
    defparam counter_4_LC_3_18_3.SEQ_MODE=4'b1010;
    defparam counter_4_LC_3_18_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_4_LC_3_18_3 (
            .in0(_gnd_net_),
            .in1(N__21770),
            .in2(_gnd_net_),
            .in3(N__21075),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(un5_counter_cry_3),
            .carryout(un5_counter_cry_4),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_5_LC_3_18_4.C_ON=1'b1;
    defparam counter_5_LC_3_18_4.SEQ_MODE=4'b1010;
    defparam counter_5_LC_3_18_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 counter_5_LC_3_18_4 (
            .in0(N__21995),
            .in1(N__21813),
            .in2(_gnd_net_),
            .in3(N__21072),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(un5_counter_cry_4),
            .carryout(un5_counter_cry_5),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_6_LC_3_18_5.C_ON=1'b1;
    defparam counter_6_LC_3_18_5.SEQ_MODE=4'b1010;
    defparam counter_6_LC_3_18_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_6_LC_3_18_5 (
            .in0(_gnd_net_),
            .in1(N__21897),
            .in2(_gnd_net_),
            .in3(N__21069),
            .lcout(counterZ0Z_6),
            .ltout(),
            .carryin(un5_counter_cry_5),
            .carryout(un5_counter_cry_6),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_7_LC_3_18_6.C_ON=1'b1;
    defparam counter_7_LC_3_18_6.SEQ_MODE=4'b1010;
    defparam counter_7_LC_3_18_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 counter_7_LC_3_18_6 (
            .in0(N__21996),
            .in1(N__21843),
            .in2(_gnd_net_),
            .in3(N__21180),
            .lcout(counterZ0Z_7),
            .ltout(),
            .carryin(un5_counter_cry_6),
            .carryout(un5_counter_cry_7),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_8_LC_3_18_7.C_ON=1'b1;
    defparam counter_8_LC_3_18_7.SEQ_MODE=4'b1010;
    defparam counter_8_LC_3_18_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 counter_8_LC_3_18_7 (
            .in0(N__21986),
            .in1(N__21855),
            .in2(_gnd_net_),
            .in3(N__21177),
            .lcout(counterZ0Z_8),
            .ltout(),
            .carryin(un5_counter_cry_7),
            .carryout(un5_counter_cry_8),
            .clk(N__46001),
            .ce(),
            .sr(N__45577));
    defparam counter_9_LC_3_19_0.C_ON=1'b1;
    defparam counter_9_LC_3_19_0.SEQ_MODE=4'b1010;
    defparam counter_9_LC_3_19_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 counter_9_LC_3_19_0 (
            .in0(N__21987),
            .in1(N__21827),
            .in2(_gnd_net_),
            .in3(N__21174),
            .lcout(counterZ0Z_9),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(un5_counter_cry_9),
            .clk(N__45993),
            .ce(),
            .sr(N__45579));
    defparam counter_10_LC_3_19_1.C_ON=1'b1;
    defparam counter_10_LC_3_19_1.SEQ_MODE=4'b1010;
    defparam counter_10_LC_3_19_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_10_LC_3_19_1 (
            .in0(_gnd_net_),
            .in1(N__21870),
            .in2(_gnd_net_),
            .in3(N__21171),
            .lcout(counterZ0Z_10),
            .ltout(),
            .carryin(un5_counter_cry_9),
            .carryout(un5_counter_cry_10),
            .clk(N__45993),
            .ce(),
            .sr(N__45579));
    defparam counter_11_LC_3_19_2.C_ON=1'b1;
    defparam counter_11_LC_3_19_2.SEQ_MODE=4'b1010;
    defparam counter_11_LC_3_19_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_11_LC_3_19_2 (
            .in0(_gnd_net_),
            .in1(N__21911),
            .in2(_gnd_net_),
            .in3(N__21168),
            .lcout(counterZ0Z_11),
            .ltout(),
            .carryin(un5_counter_cry_10),
            .carryout(un5_counter_cry_11),
            .clk(N__45993),
            .ce(),
            .sr(N__45579));
    defparam counter_12_LC_3_19_3.C_ON=1'b0;
    defparam counter_12_LC_3_19_3.SEQ_MODE=4'b1010;
    defparam counter_12_LC_3_19_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 counter_12_LC_3_19_3 (
            .in0(N__21994),
            .in1(N__21884),
            .in2(_gnd_net_),
            .in3(N__21165),
            .lcout(counterZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45993),
            .ce(),
            .sr(N__45579));
    defparam clk_10khz_LC_3_19_7.C_ON=1'b0;
    defparam clk_10khz_LC_3_19_7.SEQ_MODE=4'b1010;
    defparam clk_10khz_LC_3_19_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_10khz_LC_3_19_7 (
            .in0(_gnd_net_),
            .in1(N__21954),
            .in2(_gnd_net_),
            .in3(N__21988),
            .lcout(clk_10khz_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45993),
            .ce(),
            .sr(N__45579));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_6_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__21153),
            .in2(N__21162),
            .in3(N__23293),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_6_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__21138),
            .in2(N__21147),
            .in3(N__23314),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_6_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__21291),
            .in2(N__21303),
            .in3(N__23221),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_6_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__21276),
            .in2(N__21285),
            .in3(N__23245),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_6_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_6_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_6_4  (
            .in0(N__23269),
            .in1(N__21261),
            .in2(N__21270),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_6_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__21255),
            .in2(N__21249),
            .in3(N__23332),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_6_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__21231),
            .in2(N__21240),
            .in3(N__23173),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_6_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_6_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_6_7  (
            .in0(N__23197),
            .in1(N__21216),
            .in2(N__21225),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__21201),
            .in2(N__21210),
            .in3(N__23356),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__21186),
            .in2(N__21195),
            .in3(N__23380),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_4_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_4_7_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_4_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21354),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46068),
            .ce(),
            .sr(N__45512));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_4_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_4_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_4_8_0 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_4_8_0  (
            .in0(N__21636),
            .in1(N__23862),
            .in2(N__23622),
            .in3(N__23757),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46064),
            .ce(N__24823),
            .sr(N__45520));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_10_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_4_10_4  (
            .in0(N__21561),
            .in1(N__23794),
            .in2(_gnd_net_),
            .in3(N__23747),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46059),
            .ce(N__24775),
            .sr(N__45535));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_4_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_4_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_10_LC_4_10_5  (
            .in0(N__22911),
            .in1(N__21330),
            .in2(N__22077),
            .in3(N__21309),
            .lcout(\current_shift_inst.PI_CTRL.N_170 ),
            .ltout(\current_shift_inst.PI_CTRL.N_170_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_4_10_6 .LUT_INIT=16'b1100111011001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_4_10_6  (
            .in0(N__23588),
            .in1(N__21723),
            .in2(N__21336),
            .in3(N__23746),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46059),
            .ce(N__24775),
            .sr(N__45535));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_11_1  (
            .in0(N__22408),
            .in1(N__22446),
            .in2(N__22366),
            .in3(N__22516),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_21_LC_4_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_21_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_21_LC_4_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGGAM_21_LC_4_11_2  (
            .in0(N__22570),
            .in1(N__22230),
            .in2(N__22959),
            .in3(N__23096),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIONJC1_12_LC_4_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIONJC1_12_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIONJC1_12_LC_4_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIONJC1_12_LC_4_11_3  (
            .in0(N__21680),
            .in1(N__22473),
            .in2(N__21333),
            .in3(N__21432),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQV7U3_20_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQV7U3_20_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQV7U3_20_LC_4_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQV7U3_20_LC_4_11_4  (
            .in0(N__21324),
            .in1(N__22063),
            .in2(N__21318),
            .in3(N__23003),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_4_11_6  (
            .in0(N__22788),
            .in1(N__22622),
            .in2(N__22197),
            .in3(N__21681),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI676B_27_LC_4_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI676B_27_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI676B_27_LC_4_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI676B_27_LC_4_11_7  (
            .in0(N__22134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22680),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_4_12_0 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_4_12_0  (
            .in0(N__23688),
            .in1(N__23589),
            .in2(N__23898),
            .in3(N__21522),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(N__24774),
            .sr(N__45550));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_4_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_4_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_4_12_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_4_12_1  (
            .in0(N__21360),
            .in1(N__23844),
            .in2(_gnd_net_),
            .in3(N__23686),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(N__24774),
            .sr(N__45550));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_4_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_4_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_4_12_2 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_4_12_2  (
            .in0(N__23687),
            .in1(_gnd_net_),
            .in2(N__23897),
            .in3(N__21600),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(N__24774),
            .sr(N__45550));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_3 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_4_12_3  (
            .in0(N__21696),
            .in1(N__23843),
            .in2(N__23617),
            .in3(N__23685),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(N__24774),
            .sr(N__45550));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_4_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_4_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_4_12_4 .LUT_INIT=16'b0011001011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_4_12_4  (
            .in0(N__23690),
            .in1(N__24132),
            .in2(N__23899),
            .in3(N__21422),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(N__24774),
            .sr(N__45550));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_4_12_5 .LUT_INIT=16'b1000101010001011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_4_12_5  (
            .in0(N__21486),
            .in1(N__23851),
            .in2(N__23618),
            .in3(N__23689),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46049),
            .ce(N__24774),
            .sr(N__45550));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__21417),
            .in2(N__24131),
            .in3(N__24127),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .clk(N__46041),
            .ce(N__24821),
            .sr(N__45556));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_4_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__21377),
            .in2(N__24096),
            .in3(N__21627),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__21617),
            .in2(N__24072),
            .in3(N__21594),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__21585),
            .in2(N__24051),
            .in3(N__21552),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__21542),
            .in2(N__24030),
            .in3(N__21516),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__21506),
            .in2(N__24009),
            .in3(N__21480),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__22278),
            .in2(N__24363),
            .in3(N__21477),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__22717),
            .in2(N__24339),
            .in3(N__21474),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__23041),
            .in2(N__24315),
            .in3(N__21471),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__21462),
            .in2(N__24291),
            .in3(N__21435),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__22851),
            .in2(N__24266),
            .in3(N__21702),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__24242),
            .in2(N__22188),
            .in3(N__21699),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__22480),
            .in2(N__24222),
            .in3(N__21687),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(N__22614),
            .in2(N__24197),
            .in3(N__21684),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(N__21670),
            .in2(N__24174),
            .in3(N__21648),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(N__24548),
            .in2(N__23973),
            .in3(N__21645),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_4_15_0  (
            .in0(_gnd_net_),
            .in1(N__22773),
            .in2(N__24528),
            .in3(N__21642),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_4_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(N__22370),
            .in2(N__24498),
            .in3(N__21639),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__22415),
            .in2(N__24477),
            .in3(N__21750),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(N__22437),
            .in2(N__24453),
            .in3(N__21738),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__22992),
            .in2(N__24432),
            .in3(N__21735),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__23088),
            .in2(N__24407),
            .in3(N__21732),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(N__22509),
            .in2(N__24384),
            .in3(N__21729),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__22886),
            .in2(N__24972),
            .in3(N__21726),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__22064),
            .in2(N__24942),
            .in3(N__21711),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__22238),
            .in2(N__24916),
            .in3(N__21708),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__24905),
            .in2(N__22572),
            .in3(N__21705),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__22688),
            .in2(N__24917),
            .in3(N__21927),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__24909),
            .in2(N__22957),
            .in3(N__21924),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__22821),
            .in2(N__24918),
            .in3(N__21921),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__24913),
            .in2(N__22146),
            .in3(N__21918),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_16_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_4_16_7  (
            .in0(N__24914),
            .in1(_gnd_net_),
            .in2(N__23557),
            .in3(N__21915),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un2_counter_1_LC_4_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un2_counter_1_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un2_counter_1_LC_4_18_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \current_shift_inst.PI_CTRL.un2_counter_1_LC_4_18_0  (
            .in0(N__21912),
            .in1(N__21896),
            .in2(N__21885),
            .in3(N__22014),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un2_counterZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un2_counter_LC_4_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un2_counter_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un2_counter_LC_4_18_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un2_counter_LC_4_18_1  (
            .in0(N__21869),
            .in1(N__21801),
            .in2(N__21858),
            .in3(N__21756),
            .lcout(\current_shift_inst.PI_CTRL.un2_counterZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un2_counter_8_LC_4_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un2_counter_8_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un2_counter_8_LC_4_18_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un2_counter_8_LC_4_18_2  (
            .in0(N__21854),
            .in1(N__21842),
            .in2(N__21831),
            .in3(N__21812),
            .lcout(\current_shift_inst.PI_CTRL.un2_counterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un2_counter_7_LC_4_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un2_counter_7_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un2_counter_7_LC_4_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.un2_counter_7_LC_4_18_3  (
            .in0(N__21794),
            .in1(N__21782),
            .in2(N__21771),
            .in3(N__22033),
            .lcout(\current_shift_inst.PI_CTRL.un2_counterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1_LC_4_19_1.C_ON=1'b0;
    defparam counter_1_LC_4_19_1.SEQ_MODE=4'b1010;
    defparam counter_1_LC_4_19_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 counter_1_LC_4_19_1 (
            .in0(N__22017),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22037),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45982),
            .ce(),
            .sr(N__45578));
    defparam counter_0_LC_4_19_2.C_ON=1'b0;
    defparam counter_0_LC_4_19_2.SEQ_MODE=4'b1010;
    defparam counter_0_LC_4_19_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 counter_0_LC_4_19_2 (
            .in0(_gnd_net_),
            .in1(N__21985),
            .in2(_gnd_net_),
            .in3(N__22016),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45982),
            .ce(),
            .sr(N__45578));
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_19_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_cnv_0_LC_4_19_4  (
            .in0(N__29392),
            .in1(N__21984),
            .in2(_gnd_net_),
            .in3(N__21953),
            .lcout(N_748_g),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_4_24_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_24_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_24_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_5_6_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_5_6_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_5_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_5_6_0  (
            .in0(N__23152),
            .in1(N__23294),
            .in2(_gnd_net_),
            .in3(N__21942),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_1_LC_5_6_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_5_6_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_5_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_5_6_1  (
            .in0(N__23148),
            .in1(N__23315),
            .in2(_gnd_net_),
            .in3(N__21939),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_2_LC_5_6_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_5_6_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_5_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_5_6_2  (
            .in0(N__23153),
            .in1(N__23229),
            .in2(_gnd_net_),
            .in3(N__21936),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_3_LC_5_6_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_5_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_5_6_3  (
            .in0(N__23149),
            .in1(N__23253),
            .in2(_gnd_net_),
            .in3(N__21933),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_4_LC_5_6_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_5_6_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_5_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_5_6_4  (
            .in0(N__23154),
            .in1(N__23273),
            .in2(_gnd_net_),
            .in3(N__21930),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_5_LC_5_6_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_5_6_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_5_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_5_6_5  (
            .in0(N__23150),
            .in1(N__23336),
            .in2(_gnd_net_),
            .in3(N__22104),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_6_LC_5_6_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_5_6_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_5_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_5_6_6  (
            .in0(N__23155),
            .in1(N__23174),
            .in2(_gnd_net_),
            .in3(N__22101),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_7_LC_5_6_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_5_6_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_5_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_5_6_7  (
            .in0(N__23151),
            .in1(N__23201),
            .in2(_gnd_net_),
            .in3(N__22098),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__46069),
            .ce(),
            .sr(N__45494));
    defparam \pwm_generator_inst.counter_8_LC_5_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_5_7_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_5_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_5_7_0  (
            .in0(N__23157),
            .in1(N__23357),
            .in2(_gnd_net_),
            .in3(N__22095),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__46065),
            .ce(),
            .sr(N__45502));
    defparam \pwm_generator_inst.counter_9_LC_5_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_5_7_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_5_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_9_LC_5_7_1  (
            .in0(N__23156),
            .in1(N__23381),
            .in2(_gnd_net_),
            .in3(N__22092),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46065),
            .ce(),
            .sr(N__45502));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_5_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_5_10_5 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_5_10_5  (
            .in0(N__22089),
            .in1(N__23795),
            .in2(N__23619),
            .in3(N__23745),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46056),
            .ce(N__24871),
            .sr(N__45528));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI736M_11_LC_5_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI736M_11_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI736M_11_LC_5_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI736M_11_LC_5_11_1  (
            .in0(N__22192),
            .in1(N__23978),
            .in2(N__22623),
            .in3(N__22783),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI225B_20_LC_5_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI225B_20_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI225B_20_LC_5_11_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI225B_20_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__22056),
            .in2(_gnd_net_),
            .in3(N__22996),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_5_11_4  (
            .in0(N__22231),
            .in1(N__22138),
            .in2(N__22956),
            .in3(N__22681),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICB2E2_12_LC_5_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICB2E2_12_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICB2E2_12_LC_5_11_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICB2E2_12_LC_5_11_5  (
            .in0(N__23525),
            .in1(N__22481),
            .in2(N__22449),
            .in3(N__22323),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_5_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_5_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_5_11_6  (
            .in0(N__22445),
            .in1(N__22407),
            .in2(N__22520),
            .in3(N__22356),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQNHC1_21_LC_5_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQNHC1_21_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQNHC1_21_LC_5_11_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQNHC1_21_LC_5_11_7  (
            .in0(N__22557),
            .in1(N__23095),
            .in2(N__22332),
            .in3(N__22329),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_10_LC_5_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_10_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_10_LC_5_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_10_LC_5_12_4  (
            .in0(N__22317),
            .in1(N__22308),
            .in2(N__23943),
            .in3(N__22299),
            .lcout(\current_shift_inst.PI_CTRL.N_171 ),
            .ltout(\current_shift_inst.PI_CTRL.N_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_5_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_5_12_5 .LUT_INIT=16'b1100110001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_5_12_5  (
            .in0(N__23542),
            .in1(N__22293),
            .in2(N__22287),
            .in3(N__23863),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46042),
            .ce(N__24857),
            .sr(N__45542));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_5_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_5_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_5_13_0 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_5_13_0  (
            .in0(N__23681),
            .in1(N__23544),
            .in2(N__22257),
            .in3(N__23869),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_5_13_1 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_5_13_1  (
            .in0(N__22203),
            .in1(N__23864),
            .in2(N__23599),
            .in3(N__23678),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_5_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_5_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_5_13_3 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_5_13_3  (
            .in0(N__22158),
            .in1(N__23867),
            .in2(N__23602),
            .in3(N__23683),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_5_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_5_13_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_5_13_4  (
            .in0(N__23680),
            .in1(N__23543),
            .in2(N__22800),
            .in3(N__23868),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_5_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_5_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_5_13_5 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_5_13_5  (
            .in0(N__22752),
            .in1(N__23865),
            .in2(N__23600),
            .in3(N__23679),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_13_6 .LUT_INIT=16'b1100110000001101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_5_13_6  (
            .in0(N__23684),
            .in1(N__22746),
            .in2(N__23613),
            .in3(N__23870),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_5_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_5_13_7 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_5_13_7  (
            .in0(N__22701),
            .in1(N__23866),
            .in2(N__23601),
            .in3(N__23682),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46030),
            .ce(N__24785),
            .sr(N__45551));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_5_14_0  (
            .in0(N__24173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24243),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_5_14_2 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_5_14_2  (
            .in0(N__22629),
            .in1(N__23905),
            .in2(N__23610),
            .in3(N__23728),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_5_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_5_14_3 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_5_14_3  (
            .in0(N__23731),
            .in1(N__23565),
            .in2(N__23921),
            .in3(N__22584),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_5_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_5_14_4 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_5_14_4  (
            .in0(N__22527),
            .in1(N__23907),
            .in2(N__23612),
            .in3(N__23730),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_5_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_5_14_6 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_5_14_6  (
            .in0(N__23103),
            .in1(N__23906),
            .in2(N__23611),
            .in3(N__23729),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_5_14_7 .LUT_INIT=16'b1111001100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_5_14_7  (
            .in0(N__23732),
            .in1(N__23566),
            .in2(N__23922),
            .in3(N__23061),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46019),
            .ce(N__24856),
            .sr(N__45557));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_1 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_5_15_1  (
            .in0(N__23022),
            .in1(N__23914),
            .in2(N__23580),
            .in3(N__23733),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46011),
            .ce(N__24826),
            .sr(N__45562));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_5_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_5_15_3 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_5_15_3  (
            .in0(N__23016),
            .in1(N__23916),
            .in2(N__23582),
            .in3(N__23735),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46011),
            .ce(N__24826),
            .sr(N__45562));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_5_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_5_15_5 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_5_15_5  (
            .in0(N__23010),
            .in1(N__23915),
            .in2(N__23581),
            .in3(N__23734),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46011),
            .ce(N__24826),
            .sr(N__45562));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_5_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_5_15_6 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_5_15_6  (
            .in0(N__23736),
            .in1(N__23508),
            .in2(N__22968),
            .in3(N__23917),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46011),
            .ce(N__24826),
            .sr(N__45562));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_10_LC_5_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_10_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI99AM_10_LC_5_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI99AM_10_LC_5_16_0  (
            .in0(N__22822),
            .in1(N__22852),
            .in2(N__23524),
            .in3(N__22885),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_5_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_5_16_3 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_5_16_3  (
            .in0(N__22899),
            .in1(N__23918),
            .in2(N__23583),
            .in3(N__23755),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46002),
            .ce(N__24732),
            .sr(N__45567));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_5_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_5_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_5_16_4  (
            .in0(N__22884),
            .in1(N__22853),
            .in2(N__22829),
            .in3(N__23974),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_5 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_5_16_5  (
            .in0(N__23928),
            .in1(N__23919),
            .in2(N__23584),
            .in3(N__23756),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46002),
            .ce(N__24732),
            .sr(N__45567));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_7_4_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_7_4_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_7_4_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23397),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46070),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_7_6_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_7_6_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNITBL3_9_LC_7_6_0  (
            .in0(N__23385),
            .in1(N__23361),
            .in2(_gnd_net_),
            .in3(N__23337),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_7_6_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_7_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIRPD2_0_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__23316),
            .in2(_gnd_net_),
            .in3(N__23295),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_7_6_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_7_6_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_2_LC_7_6_2  (
            .in0(N__23274),
            .in1(N__23252),
            .in2(N__23232),
            .in3(N__23228),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_7_6_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_7_6_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_6_LC_7_6_3  (
            .in0(N__23208),
            .in1(N__23202),
            .in2(N__23181),
            .in3(N__23178),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_7_11_0  (
            .in0(N__29038),
            .in1(N__28822),
            .in2(N__25104),
            .in3(N__28964),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46031),
            .ce(),
            .sr(N__45521));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_7_11_2  (
            .in0(N__29037),
            .in1(N__28821),
            .in2(_gnd_net_),
            .in3(N__28963),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_tr.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_7_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_7_11_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_7_11_3  (
            .in0(N__25016),
            .in1(N__29193),
            .in2(N__24153),
            .in3(N__29158),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46031),
            .ce(),
            .sr(N__45521));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24068),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46020),
            .ce(N__24846),
            .sr(N__45529));
    defparam \current_shift_inst.control_input_0_LC_7_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_0_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_0_LC_7_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_0_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__25185),
            .in2(N__26970),
            .in3(N__26969),
            .lcout(\current_shift_inst.control_inputZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\current_shift_inst.control_input_1_cry_0 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_1_LC_7_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_1_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_1_LC_7_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_1_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__25260),
            .in2(_gnd_net_),
            .in3(N__24075),
            .lcout(\current_shift_inst.control_inputZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_0 ),
            .carryout(\current_shift_inst.control_input_1_cry_1 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_2_LC_7_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_2_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_2_LC_7_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_2_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__25155),
            .in2(_gnd_net_),
            .in3(N__24054),
            .lcout(\current_shift_inst.control_inputZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_1 ),
            .carryout(\current_shift_inst.control_input_1_cry_2 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_3_LC_7_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_3_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_3_LC_7_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_3_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__25173),
            .in2(_gnd_net_),
            .in3(N__24033),
            .lcout(\current_shift_inst.control_inputZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_2 ),
            .carryout(\current_shift_inst.control_input_1_cry_3 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_4_LC_7_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_4_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_4_LC_7_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_4_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__25239),
            .in2(_gnd_net_),
            .in3(N__24012),
            .lcout(\current_shift_inst.control_inputZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_3 ),
            .carryout(\current_shift_inst.control_input_1_cry_4 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_5_LC_7_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_5_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_5_LC_7_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_5_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__25143),
            .in2(_gnd_net_),
            .in3(N__23988),
            .lcout(\current_shift_inst.control_inputZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_4 ),
            .carryout(\current_shift_inst.control_input_1_cry_5 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_6_LC_7_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_6_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_6_LC_7_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_6_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__25149),
            .in2(_gnd_net_),
            .in3(N__24342),
            .lcout(\current_shift_inst.control_inputZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_5 ),
            .carryout(\current_shift_inst.control_input_1_cry_6 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_7_LC_7_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_7_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_7_LC_7_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_7_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__25227),
            .in2(_gnd_net_),
            .in3(N__24318),
            .lcout(\current_shift_inst.control_inputZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_6 ),
            .carryout(\current_shift_inst.control_input_1_cry_7 ),
            .clk(N__46012),
            .ce(N__24825),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_8_LC_7_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_8_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_8_LC_7_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_8_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__25200),
            .in2(_gnd_net_),
            .in3(N__24294),
            .lcout(\current_shift_inst.control_inputZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\current_shift_inst.control_input_1_cry_8 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_9_LC_7_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_9_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_9_LC_7_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_9_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__25272),
            .in2(_gnd_net_),
            .in3(N__24270),
            .lcout(\current_shift_inst.control_inputZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_8 ),
            .carryout(\current_shift_inst.control_input_1_cry_9 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_10_LC_7_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_10_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_10_LC_7_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_10_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__25113),
            .in2(_gnd_net_),
            .in3(N__24246),
            .lcout(\current_shift_inst.control_inputZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_9 ),
            .carryout(\current_shift_inst.control_input_1_cry_10 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_11_LC_7_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_11_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_11_LC_7_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.control_input_11_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25209),
            .in3(N__24225),
            .lcout(\current_shift_inst.control_inputZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_10 ),
            .carryout(\current_shift_inst.control_input_1_cry_11 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_12_LC_7_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_12_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_12_LC_7_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_12_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__25125),
            .in2(_gnd_net_),
            .in3(N__24201),
            .lcout(\current_shift_inst.control_inputZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_11 ),
            .carryout(\current_shift_inst.control_input_1_cry_12 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_13_LC_7_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_13_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_13_LC_7_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_13_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__25131),
            .in2(_gnd_net_),
            .in3(N__24177),
            .lcout(\current_shift_inst.control_inputZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_12 ),
            .carryout(\current_shift_inst.control_input_1_cry_13 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_14_LC_7_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_14_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_14_LC_7_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_14_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__25137),
            .in2(_gnd_net_),
            .in3(N__24156),
            .lcout(\current_shift_inst.control_inputZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_13 ),
            .carryout(\current_shift_inst.control_input_1_cry_14 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_15_LC_7_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_15_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_15_LC_7_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_15_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__25119),
            .in2(_gnd_net_),
            .in3(N__24531),
            .lcout(\current_shift_inst.control_inputZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_14 ),
            .carryout(\current_shift_inst.control_input_1_cry_15 ),
            .clk(N__46003),
            .ce(N__24845),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_16_LC_7_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_16_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_16_LC_7_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_16_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__25215),
            .in2(_gnd_net_),
            .in3(N__24501),
            .lcout(\current_shift_inst.control_inputZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\current_shift_inst.control_input_1_cry_16 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_17_LC_7_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_17_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_17_LC_7_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_17_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__25248),
            .in2(_gnd_net_),
            .in3(N__24480),
            .lcout(\current_shift_inst.control_inputZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_16 ),
            .carryout(\current_shift_inst.control_input_1_cry_17 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_18_LC_7_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_18_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_18_LC_7_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_18_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__25296),
            .in2(_gnd_net_),
            .in3(N__24456),
            .lcout(\current_shift_inst.control_inputZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_17 ),
            .carryout(\current_shift_inst.control_input_1_cry_18 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_19_LC_7_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_19_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_19_LC_7_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_19_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__25287),
            .in2(_gnd_net_),
            .in3(N__24435),
            .lcout(\current_shift_inst.control_inputZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_18 ),
            .carryout(\current_shift_inst.control_input_1_cry_19 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_20_LC_7_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_20_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_20_LC_7_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_20_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__25194),
            .in2(_gnd_net_),
            .in3(N__24411),
            .lcout(\current_shift_inst.control_inputZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_19 ),
            .carryout(\current_shift_inst.control_input_1_cry_20 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_21_LC_7_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_21_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_21_LC_7_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_21_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__25059),
            .in2(_gnd_net_),
            .in3(N__24387),
            .lcout(\current_shift_inst.control_inputZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_20 ),
            .carryout(\current_shift_inst.control_input_1_cry_21 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_22_LC_7_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_22_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_22_LC_7_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_22_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(N__25065),
            .in2(_gnd_net_),
            .in3(N__24366),
            .lcout(\current_shift_inst.control_inputZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_21 ),
            .carryout(\current_shift_inst.control_input_1_cry_22 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_23_LC_7_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_23_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_23_LC_7_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_23_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__24585),
            .in2(_gnd_net_),
            .in3(N__24945),
            .lcout(\current_shift_inst.control_inputZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_1_cry_22 ),
            .carryout(\current_shift_inst.control_input_1_cry_23 ),
            .clk(N__45994),
            .ce(N__24861),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_24_LC_7_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.control_input_24_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_24_LC_7_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.control_input_24_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__25278),
            .in2(_gnd_net_),
            .in3(N__24924),
            .lcout(\current_shift_inst.control_inputZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\current_shift_inst.control_input_1_cry_24 ),
            .clk(N__45983),
            .ce(N__24805),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_25_LC_7_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_25_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \current_shift_inst.control_input_25_LC_7_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.control_input_25_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__25626),
            .in2(_gnd_net_),
            .in3(N__24921),
            .lcout(\current_shift_inst.control_inputZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45983),
            .ce(N__24805),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_7_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_7_17_4 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_7_17_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__29383),
            .in2(_gnd_net_),
            .in3(N__38186),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45976),
            .ce(),
            .sr(N__45563));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_7_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_7_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_7_18_2  (
            .in0(N__29814),
            .in1(N__32292),
            .in2(N__30333),
            .in3(N__27807),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_7_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_7_20_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_7_20_2  (
            .in0(N__29802),
            .in1(N__32526),
            .in2(N__30334),
            .in3(N__27897),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_22_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_7_22_6  (
            .in0(N__25650),
            .in1(N__26187),
            .in2(_gnd_net_),
            .in3(N__27092),
            .lcout(\current_shift_inst.control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24573),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46062),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_7_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_7_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24564),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46057),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_8_9_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_8_9_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_8_9_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_8_9_2 (
            .in0(N__25026),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46043),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_8_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_8_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__25017),
            .in2(_gnd_net_),
            .in3(N__24995),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_8_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_8_10_0 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_8_10_0  (
            .in0(N__27497),
            .in1(N__29059),
            .in2(N__25167),
            .in3(N__38213),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46032),
            .ce(),
            .sr(N__45503));
    defparam \phase_controller_inst2.state_0_LC_8_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_8_10_4 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst2.state_0_LC_8_10_4  (
            .in0(N__31792),
            .in1(N__25015),
            .in2(N__31739),
            .in3(N__24996),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46032),
            .ce(),
            .sr(N__45503));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__25074),
            .in2(N__26316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_8_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_8_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__26289),
            .in2(_gnd_net_),
            .in3(N__24984),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_8_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_3_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__25083),
            .in2(N__26271),
            .in3(N__24981),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_8_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_8_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_4_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__26250),
            .in2(_gnd_net_),
            .in3(N__24978),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_8_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_8_11_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_5_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26499),
            .in3(N__24975),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_8_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_8_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_6_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__26478),
            .in2(_gnd_net_),
            .in3(N__25053),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_8_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_8_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_7_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__26460),
            .in2(_gnd_net_),
            .in3(N__25050),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_8_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_8_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_8_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__26433),
            .in2(_gnd_net_),
            .in3(N__25047),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_8_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_8_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_9_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__26403),
            .in2(_gnd_net_),
            .in3(N__25044),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_9 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_8_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_8_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_10_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__26385),
            .in2(_gnd_net_),
            .in3(N__25041),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_8_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_8_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_11_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__26352),
            .in2(_gnd_net_),
            .in3(N__25038),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_8_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_8_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_12_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__26334),
            .in2(_gnd_net_),
            .in3(N__25035),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_8_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_8_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_13_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__26655),
            .in2(_gnd_net_),
            .in3(N__25032),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_8_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_8_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_14_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__26637),
            .in2(_gnd_net_),
            .in3(N__25029),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_8_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_8_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_15_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(N__26619),
            .in2(_gnd_net_),
            .in3(N__25107),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_8_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_8_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_16_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(N__26585),
            .in2(_gnd_net_),
            .in3(N__25095),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_8_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_17_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__26565),
            .in2(_gnd_net_),
            .in3(N__25092),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_17 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_8_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_18_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__26547),
            .in2(_gnd_net_),
            .in3(N__25089),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_8_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_8_13_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_19_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__26529),
            .in2(_gnd_net_),
            .in3(N__25086),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJ_LC_8_13_5  (
            .in0(N__29182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29148),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_RNIF9HJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_13_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_8_13_7  (
            .in0(N__29181),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29147),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_14_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_8_14_0  (
            .in0(N__27083),
            .in1(N__26202),
            .in2(_gnd_net_),
            .in3(N__25668),
            .lcout(\current_shift_inst.control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_14_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_8_14_1  (
            .in0(N__25680),
            .in1(N__26217),
            .in2(_gnd_net_),
            .in3(N__27082),
            .lcout(\current_shift_inst.control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_8_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_8_14_3 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_8_14_3  (
            .in0(N__25992),
            .in1(N__25455),
            .in2(_gnd_net_),
            .in3(N__27079),
            .lcout(\current_shift_inst.control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_14_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__31722),
            .in2(_gnd_net_),
            .in3(N__31793),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_8_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_8_14_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_8_14_5  (
            .in0(N__25311),
            .in1(N__25851),
            .in2(_gnd_net_),
            .in3(N__27078),
            .lcout(\current_shift_inst.control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_8_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_8_14_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_8_14_6  (
            .in0(N__27081),
            .in1(N__25950),
            .in2(_gnd_net_),
            .in3(N__25419),
            .lcout(\current_shift_inst.control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_8_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_8_14_7 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_8_14_7  (
            .in0(N__25965),
            .in1(N__25431),
            .in2(_gnd_net_),
            .in3(N__27080),
            .lcout(\current_shift_inst.control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_15_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_8_15_0  (
            .in0(N__27089),
            .in1(N__25539),
            .in2(_gnd_net_),
            .in3(N__26091),
            .lcout(\current_shift_inst.control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_8_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_8_15_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_8_15_1  (
            .in0(N__26109),
            .in1(N__25551),
            .in2(_gnd_net_),
            .in3(N__27088),
            .lcout(\current_shift_inst.control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_8_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_8_15_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_8_15_2  (
            .in0(N__27087),
            .in1(N__26124),
            .in2(_gnd_net_),
            .in3(N__25566),
            .lcout(\current_shift_inst.control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_15_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_8_15_3  (
            .in0(N__25527),
            .in1(N__26076),
            .in2(_gnd_net_),
            .in3(N__27090),
            .lcout(\current_shift_inst.control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_8_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_8_15_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_8_15_4  (
            .in0(N__27085),
            .in1(N__25368),
            .in2(_gnd_net_),
            .in3(N__25890),
            .lcout(\current_shift_inst.control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_8_15_5  (
            .in0(N__25512),
            .in1(N__26061),
            .in2(_gnd_net_),
            .in3(N__27091),
            .lcout(\current_shift_inst.control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_8_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_8_15_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_8_15_6  (
            .in0(N__27086),
            .in1(N__26139),
            .in2(_gnd_net_),
            .in3(N__25587),
            .lcout(\current_shift_inst.control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_8_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_8_15_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_8_15_7  (
            .in0(N__25395),
            .in1(N__25923),
            .in2(_gnd_net_),
            .in3(N__27084),
            .lcout(\current_shift_inst.control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_8_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_8_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32511),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_8_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_8_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_8_16_4  (
            .in0(N__29591),
            .in1(N__31566),
            .in2(N__30493),
            .in3(N__30729),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_16_5 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_8_16_5  (
            .in0(N__26232),
            .in1(N__25704),
            .in2(_gnd_net_),
            .in3(N__27077),
            .lcout(\current_shift_inst.control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_8_16_6 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_8_16_6  (
            .in0(N__32484),
            .in1(N__30332),
            .in2(N__29696),
            .in3(N__27867),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_8_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_8_17_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_8_17_0  (
            .in0(N__25875),
            .in1(N__25338),
            .in2(_gnd_net_),
            .in3(N__27018),
            .lcout(\current_shift_inst.control_input_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_8_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_8_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_8_17_1  (
            .in0(N__29801),
            .in1(N__32757),
            .in2(N__30492),
            .in3(N__27978),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_8_17_3  (
            .in0(N__27020),
            .in1(N__26031),
            .in2(_gnd_net_),
            .in3(N__25482),
            .lcout(\current_shift_inst.control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_8_17_4  (
            .in0(N__26016),
            .in1(N__25467),
            .in2(_gnd_net_),
            .in3(N__27021),
            .lcout(\current_shift_inst.control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_8_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_8_17_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNI9GMC2_LC_8_17_5  (
            .in0(N__27022),
            .in1(N__25641),
            .in2(_gnd_net_),
            .in3(N__26175),
            .lcout(\current_shift_inst.control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_8_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_8_17_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_8_17_6  (
            .in0(N__25380),
            .in1(N__25905),
            .in2(_gnd_net_),
            .in3(N__27019),
            .lcout(\current_shift_inst.control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_8_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_8_18_3 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_8_18_3  (
            .in0(N__25860),
            .in1(N__25320),
            .in2(_gnd_net_),
            .in3(N__27023),
            .lcout(\current_shift_inst.control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_8_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_8_18_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_8_18_4  (
            .in0(N__27026),
            .in1(N__25494),
            .in2(_gnd_net_),
            .in3(N__26046),
            .lcout(\current_shift_inst.control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_18_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_8_18_5  (
            .in0(N__25443),
            .in1(N__25977),
            .in2(_gnd_net_),
            .in3(N__27024),
            .lcout(\current_shift_inst.control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_8_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_8_18_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_8_18_6  (
            .in0(N__27025),
            .in1(N__25935),
            .in2(_gnd_net_),
            .in3(N__25407),
            .lcout(\current_shift_inst.control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_8_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_8_18_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_8_18_7  (
            .in0(N__29692),
            .in1(N__27633),
            .in2(N__26762),
            .in3(N__26703),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__27528),
            .in2(N__34179),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__25353),
            .in2(N__26755),
            .in3(N__34618),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_19_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_19_2  (
            .in0(N__34619),
            .in1(N__29235),
            .in2(N__30348),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_8_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__30145),
            .in2(N__26943),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_8_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__28413),
            .in2(N__30349),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_8_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__25347),
            .in2(N__30272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__26835),
            .in2(N__30350),
            .in3(N__25329),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__25326),
            .in2(N__30273),
            .in3(N__25314),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__27249),
            .in2(N__30278),
            .in3(N__25299),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__26871),
            .in2(N__30282),
            .in3(N__25446),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__28350),
            .in2(N__30279),
            .in3(N__25434),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__28317),
            .in2(N__30283),
            .in3(N__25422),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__26910),
            .in2(N__30280),
            .in3(N__25410),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__27240),
            .in2(N__30284),
            .in3(N__25398),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__28281),
            .in2(N__30281),
            .in3(N__25383),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_20_7  (
            .in0(_gnd_net_),
            .in1(N__28245),
            .in2(N__30285),
            .in3(N__25371),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(N__28566),
            .in2(N__30464),
            .in3(N__25356),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(N__25593),
            .in2(N__30438),
            .in3(N__25578),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(N__25575),
            .in2(N__30465),
            .in3(N__25554),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(N__28062),
            .in2(N__30439),
            .in3(N__25542),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_21_4  (
            .in0(_gnd_net_),
            .in1(N__28098),
            .in2(N__30466),
            .in3(N__25530),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_21_5  (
            .in0(_gnd_net_),
            .in1(N__28449),
            .in2(N__30440),
            .in3(N__25515),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_21_6  (
            .in0(_gnd_net_),
            .in1(N__27306),
            .in2(N__30467),
            .in3(N__25497),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(N__28026),
            .in2(N__30441),
            .in3(N__25485),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(N__28188),
            .in2(N__30595),
            .in3(N__25470),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(N__30448),
            .in2(N__27213),
            .in3(N__25707),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__28158),
            .in2(N__30596),
            .in3(N__25692),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(N__25689),
            .in2(N__30468),
            .in3(N__25671),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(N__28386),
            .in2(N__30597),
            .in3(N__25653),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(N__27297),
            .in2(N__30469),
            .in3(N__25644),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_8_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_8_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_8_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNII18T_LC_8_22_6  (
            .in0(_gnd_net_),
            .in1(N__28545),
            .in2(N__30598),
            .in3(N__25632),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_0_25_LC_8_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_8_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_0_25_LC_8_22_7 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \current_shift_inst.control_input_RNO_0_25_LC_8_22_7  (
            .in0(N__27681),
            .in1(N__27093),
            .in2(N__26157),
            .in3(N__25629),
            .lcout(\current_shift_inst.control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_8_29_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_8_29_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_8_29_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_8_29_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31743),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45930),
            .ce(),
            .sr(N__45581));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_9_7_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_9_7_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_9_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_9_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25602),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46050),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_9_7_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_9_7_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_9_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25761),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46050),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_9_10_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_9_10_0  (
            .in0(N__28824),
            .in1(N__28944),
            .in2(N__29084),
            .in3(N__25749),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(),
            .sr(N__45495));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_9_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_9_10_1 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_9_10_1  (
            .in0(N__28942),
            .in1(N__29039),
            .in2(N__25743),
            .in3(N__28825),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(),
            .sr(N__45495));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_9_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_9_10_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_9_10_2  (
            .in0(N__28823),
            .in1(N__28943),
            .in2(N__29083),
            .in3(N__25734),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46021),
            .ce(),
            .sr(N__45495));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_9_11_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_9_11_0  (
            .in0(N__28814),
            .in1(N__28935),
            .in2(N__29085),
            .in3(N__25728),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_9_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_RNO_0_1_LC_9_11_1  (
            .in0(N__29189),
            .in1(N__26315),
            .in2(_gnd_net_),
            .in3(N__29152),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_9_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_9_11_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_9_11_2  (
            .in0(N__28817),
            .in1(N__29058),
            .in2(N__25722),
            .in3(N__28941),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_9_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_9_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_9_11_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_9_11_3  (
            .in0(N__25719),
            .in1(N__29046),
            .in2(N__28965),
            .in3(N__28820),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_9_11_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_9_11_4  (
            .in0(N__28815),
            .in1(N__28936),
            .in2(N__29086),
            .in3(N__25713),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_9_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_9_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_9_11_5 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_9_11_5  (
            .in0(N__28933),
            .in1(N__29047),
            .in2(N__25821),
            .in3(N__28818),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_9_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_9_11_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_9_11_6  (
            .in0(N__28816),
            .in1(N__28937),
            .in2(N__29087),
            .in3(N__25812),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_9_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_9_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_9_11_7 .LUT_INIT=16'b1110000010110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_9_11_7  (
            .in0(N__28934),
            .in1(N__29048),
            .in2(N__25806),
            .in3(N__28819),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46013),
            .ce(),
            .sr(N__45504));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_9_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_9_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_9_12_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_9_12_0  (
            .in0(N__28826),
            .in1(N__29099),
            .in2(N__28978),
            .in3(N__25797),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_9_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_9_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_9_12_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_9_12_1  (
            .in0(N__28945),
            .in1(N__28830),
            .in2(N__29110),
            .in3(N__25791),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_9_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_9_12_2 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_9_12_2  (
            .in0(N__28827),
            .in1(N__29100),
            .in2(N__28979),
            .in3(N__25785),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_9_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_9_12_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_9_12_3  (
            .in0(N__25779),
            .in1(N__28831),
            .in2(N__28967),
            .in3(N__29094),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_9_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_9_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_9_12_4 .LUT_INIT=16'b1010100010001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_9_12_4  (
            .in0(N__25773),
            .in1(N__28946),
            .in2(N__28836),
            .in3(N__29101),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_9_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_9_12_5 .LUT_INIT=16'b1100100011000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_9_12_5  (
            .in0(N__29103),
            .in1(N__25767),
            .in2(N__28968),
            .in3(N__28832),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_9_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_9_12_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_9_12_6  (
            .in0(N__28828),
            .in1(N__29102),
            .in2(N__28980),
            .in3(N__25833),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_9_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_9_12_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_9_12_7  (
            .in0(N__29098),
            .in1(N__28829),
            .in2(N__28966),
            .in3(N__25827),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46004),
            .ce(),
            .sr(N__45513));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_13_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_13_2  (
            .in0(N__29579),
            .in1(N__32204),
            .in2(N__30672),
            .in3(N__27771),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_13_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__32994),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45995),
            .ce(N__32967),
            .sr(N__45522));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_9_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33666),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45984),
            .ce(N__32966),
            .sr(N__45530));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__34652),
            .in2(N__34623),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__26679),
            .in2(N__34580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__26673),
            .in2(N__34588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__26847),
            .in2(N__34581),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__26811),
            .in2(N__34589),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__26859),
            .in2(N__34582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__26775),
            .in2(N__34590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__26709),
            .in2(N__34583),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__26841),
            .in2(N__34579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__26817),
            .in2(N__34587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__26928),
            .in2(N__34576),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__26853),
            .in2(N__34584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__26823),
            .in2(N__34577),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__26922),
            .in2(N__34585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__26898),
            .in2(N__34578),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(N__26916),
            .in2(N__34586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__26877),
            .in2(N__34567),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__26892),
            .in2(N__34571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__27135),
            .in2(N__34568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__34490),
            .in2(N__26886),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__27129),
            .in2(N__34569),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__30807),
            .in2(N__34572),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__27123),
            .in2(N__34570),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__27117),
            .in2(N__34573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__34375),
            .in2(N__27144),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__27111),
            .in2(N__34478),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__28131),
            .in2(N__34481),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__26949),
            .in2(N__34479),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__27219),
            .in2(N__34482),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__27174),
            .in2(N__34480),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__28224),
            .in2(N__34483),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__29767),
            .in2(_gnd_net_),
            .in3(N__25836),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__34206),
            .in2(N__34178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__26721),
            .in2(N__26754),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__27159),
            .in2(N__30346),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_9_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__27279),
            .in2(N__30424),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_9_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__30186),
            .in2(N__27168),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_9_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__30705),
            .in2(N__30425),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__29448),
            .in2(N__30347),
            .in3(N__25863),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__30141),
            .in2(N__27153),
            .in3(N__25854),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__28461),
            .in2(N__30274),
            .in3(N__25839),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__26001),
            .in2(N__30426),
            .in3(N__25980),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__27273),
            .in2(N__30275),
            .in3(N__25968),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__27336),
            .in2(N__30427),
            .in3(N__25953),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__27348),
            .in2(N__30276),
            .in3(N__25938),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__27267),
            .in2(N__30428),
            .in3(N__25926),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__27285),
            .in2(N__30277),
            .in3(N__25908),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__27354),
            .in2(N__30429),
            .in3(N__25893),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__28236),
            .in2(N__30430),
            .in3(N__25878),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__27255),
            .in2(N__30434),
            .in3(N__26127),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__27105),
            .in2(N__30431),
            .in3(N__26112),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__27318),
            .in2(N__30435),
            .in3(N__26094),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__27342),
            .in2(N__30432),
            .in3(N__26079),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__27330),
            .in2(N__30436),
            .in3(N__26064),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__27312),
            .in2(N__30433),
            .in3(N__26049),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__27261),
            .in2(N__30437),
            .in3(N__26034),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(N__30238),
            .in2(N__27513),
            .in3(N__26019),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__27198),
            .in2(N__30442),
            .in3(N__26004),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__28176),
            .in2(N__30458),
            .in3(N__26220),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__27186),
            .in2(N__30443),
            .in3(N__26205),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__27231),
            .in2(N__30459),
            .in3(N__26190),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__27324),
            .in2(N__30444),
            .in3(N__26178),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_9_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_9_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIJ39T_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__28544),
            .in2(N__30460),
            .in3(N__26163),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_2_25_LC_9_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_2_25_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_2_25_LC_9_22_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.control_input_RNO_2_25_LC_9_22_7  (
            .in0(N__29809),
            .in1(N__30268),
            .in2(_gnd_net_),
            .in3(N__26160),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_27_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27486),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45932),
            .ce(),
            .sr(N__45580));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_10_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__31464),
            .in2(_gnd_net_),
            .in3(N__33258),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46014),
            .ce(N__29322),
            .sr(N__45480));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_10_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_10_10_0  (
            .in0(N__31463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33327),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46006),
            .ce(N__29321),
            .sr(N__45485));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_10_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__31886),
            .in2(_gnd_net_),
            .in3(N__35841),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46006),
            .ce(N__29321),
            .sr(N__45485));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_10_4 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_10_10_4  (
            .in0(N__28704),
            .in1(N__35949),
            .in2(N__31895),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46006),
            .ce(N__29321),
            .sr(N__45485));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_10_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_10_10_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_10_10_6  (
            .in0(N__31890),
            .in1(N__35907),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46006),
            .ce(N__29321),
            .sr(N__45485));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_10_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_10_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38076),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46006),
            .ce(N__29321),
            .sr(N__45485));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_10_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_10_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_10_11_0  (
            .in0(_gnd_net_),
            .in1(N__26295),
            .in2(N__27384),
            .in3(N__26311),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_10_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_10_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(N__26277),
            .in2(N__27393),
            .in3(N__26288),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_10_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_10_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__26256),
            .in2(N__27552),
            .in3(N__26267),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_10_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_10_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(N__26238),
            .in2(N__27366),
            .in3(N__26249),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_10_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_10_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__26484),
            .in2(N__26511),
            .in3(N__26495),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_10_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_10_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(N__26466),
            .in2(N__27582),
            .in3(N__26477),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_10_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_10_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_10_11_6  (
            .in0(N__26459),
            .in1(N__26439),
            .in2(N__26448),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_10_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_10_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_10_11_7  (
            .in0(N__26432),
            .in1(N__26409),
            .in2(N__26421),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_10_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_10_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__26391),
            .in2(N__27375),
            .in3(N__26402),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_10_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_10_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__26373),
            .in2(N__27564),
            .in3(N__26384),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_10_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_10_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__26340),
            .in2(N__26367),
            .in3(N__26351),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_10_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_10_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__26322),
            .in2(N__27573),
            .in3(N__26333),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_10_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_10_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__26643),
            .in2(N__26667),
            .in3(N__26654),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_10_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_10_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__26625),
            .in2(N__27408),
            .in3(N__26636),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_10_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_10_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__26607),
            .in2(N__27543),
            .in3(N__26618),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_10_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_10_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(N__26571),
            .in2(N__26601),
            .in3(N__26589),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_10_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_10_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_10_13_0  (
            .in0(N__26564),
            .in1(N__26553),
            .in2(N__26802),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_10_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_10_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_10_13_1  (
            .in0(N__26546),
            .in1(N__26535),
            .in2(N__26793),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_10_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_10_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__26517),
            .in2(N__26784),
            .in3(N__26528),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26805),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_10_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43775),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45977),
            .ce(N__29316),
            .sr(N__45505));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_10_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43557),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45977),
            .ce(N__29316),
            .sr(N__45505));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_10_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38043),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45977),
            .ce(N__29316),
            .sr(N__45505));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__26694),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_14_1  (
            .in0(N__30910),
            .in1(N__32332),
            .in2(_gnd_net_),
            .in3(N__29464),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_14_2 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_10_14_2  (
            .in0(N__27626),
            .in1(N__26696),
            .in2(N__26769),
            .in3(N__29534),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_10_14_3  (
            .in0(N__30911),
            .in1(N__32287),
            .in2(_gnd_net_),
            .in3(N__27793),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_14_4 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_10_14_4  (
            .in0(N__27625),
            .in1(N__26695),
            .in2(_gnd_net_),
            .in3(N__30907),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_14_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_14_5  (
            .in0(N__30908),
            .in1(N__31679),
            .in2(_gnd_net_),
            .in3(N__29251),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_10_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_10_14_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_10_14_6  (
            .in0(N__30673),
            .in1(N__29535),
            .in2(N__32208),
            .in3(N__27764),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_14_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_14_7  (
            .in0(N__30909),
            .in1(N__31562),
            .in2(_gnd_net_),
            .in3(N__30721),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_15_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_10_15_0  (
            .in0(N__32119),
            .in1(N__30918),
            .in2(_gnd_net_),
            .in3(N__28330),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_1 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_10_15_1  (
            .in0(N__31633),
            .in1(_gnd_net_),
            .in2(N__30942),
            .in3(N__27601),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_15_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_15_2  (
            .in0(N__32236),
            .in1(N__30916),
            .in2(_gnd_net_),
            .in3(N__28474),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_15_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_10_15_3  (
            .in0(N__30494),
            .in1(N__29732),
            .in2(N__32337),
            .in3(N__29465),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_15_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_10_15_4  (
            .in0(N__32084),
            .in1(N__30919),
            .in2(_gnd_net_),
            .in3(N__27730),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_10_15_5  (
            .in0(N__30917),
            .in1(N__32197),
            .in2(_gnd_net_),
            .in3(N__27763),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_10_15_6  (
            .in0(N__31600),
            .in1(N__30915),
            .in2(_gnd_net_),
            .in3(N__28426),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_10_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_10_15_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_10_15_7  (
            .in0(N__31634),
            .in1(N__29731),
            .in2(N__30610),
            .in3(N__27602),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_0 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_16_0  (
            .in0(N__32167),
            .in1(N__28363),
            .in2(_gnd_net_),
            .in3(N__30920),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_16_1  (
            .in0(N__30921),
            .in1(N__32041),
            .in2(_gnd_net_),
            .in3(N__27695),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_10_16_2  (
            .in0(N__32605),
            .in1(N__30923),
            .in2(_gnd_net_),
            .in3(N__28261),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_10_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_10_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_10_16_3  (
            .in0(N__29630),
            .in1(N__32080),
            .in2(N__30692),
            .in3(N__27731),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_16_4  (
            .in0(N__32644),
            .in1(N__30922),
            .in2(_gnd_net_),
            .in3(N__28297),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_16_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_10_16_5  (
            .in0(N__30925),
            .in1(N__32521),
            .in2(_gnd_net_),
            .in3(N__27881),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_10_16_6  (
            .in0(N__32446),
            .in1(N__30926),
            .in2(_gnd_net_),
            .in3(N__28075),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_16_7  (
            .in0(N__30924),
            .in1(N__32568),
            .in2(_gnd_net_),
            .in3(N__28577),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_17_0  (
            .in0(N__30947),
            .in1(N__32867),
            .in2(_gnd_net_),
            .in3(N__28204),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_10_17_1  (
            .in0(N__30943),
            .in1(N__32473),
            .in2(_gnd_net_),
            .in3(N__27862),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_17_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_17_2  (
            .in0(N__30945),
            .in1(N__32404),
            .in2(_gnd_net_),
            .in3(N__28111),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3  (
            .in0(N__32932),
            .in1(N__30946),
            .in2(_gnd_net_),
            .in3(N__27827),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_17_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_10_17_4  (
            .in0(N__32899),
            .in1(N__30944),
            .in2(_gnd_net_),
            .in3(N__28039),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_10_17_5  (
            .in0(N__29697),
            .in1(N__32818),
            .in2(_gnd_net_),
            .in3(N__27997),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_17_6 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_17_6  (
            .in0(N__27863),
            .in1(N__29698),
            .in2(N__32480),
            .in3(N__30679),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27017),
            .lcout(\current_shift_inst.N_1819_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_0  (
            .in0(N__29733),
            .in1(N__32749),
            .in2(_gnd_net_),
            .in3(N__27973),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_18_1 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_18_1  (
            .in0(N__28400),
            .in1(N__29736),
            .in2(N__32723),
            .in3(N__30471),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_10_18_2  (
            .in0(N__29734),
            .in1(N__32716),
            .in2(_gnd_net_),
            .in3(N__28399),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_3  (
            .in0(N__29705),
            .in1(N__27998),
            .in2(N__30602),
            .in3(N__32819),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_18_4 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_18_4  (
            .in0(N__27999),
            .in1(N__29706),
            .in2(N__32823),
            .in3(N__30475),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_18_5 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_18_5  (
            .in0(N__27974),
            .in1(N__29735),
            .in2(N__32756),
            .in3(N__30470),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_10_18_6  (
            .in0(N__32680),
            .in1(N__29704),
            .in2(_gnd_net_),
            .in3(N__27943),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_10_18_7  (
            .in0(N__29703),
            .in1(N__31608),
            .in2(N__30603),
            .in3(N__28437),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_19_1  (
            .in0(N__29699),
            .in1(N__31680),
            .in2(N__30624),
            .in3(N__29259),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_19_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_19_2  (
            .in0(N__29707),
            .in1(N__32291),
            .in2(N__30620),
            .in3(N__27806),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_19_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_19_3  (
            .in0(N__27950),
            .in1(N__29709),
            .in2(N__30623),
            .in3(N__32688),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_4  (
            .in0(N__32646),
            .in1(N__29702),
            .in2(N__30621),
            .in3(N__28308),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_19_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_10_19_5  (
            .in0(N__29700),
            .in1(N__31641),
            .in2(N__30625),
            .in3(N__27609),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_19_6  (
            .in0(N__29708),
            .in1(N__32169),
            .in2(N__30619),
            .in3(N__28374),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_19_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_10_19_7  (
            .in0(N__29701),
            .in1(N__32045),
            .in2(N__30622),
            .in3(N__27707),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_20_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_20_0  (
            .in0(N__29821),
            .in1(N__32906),
            .in2(N__30678),
            .in3(N__28050),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_20_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_20_1  (
            .in0(N__32522),
            .in1(N__29820),
            .in2(N__30667),
            .in3(N__27893),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_20_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_10_20_3  (
            .in0(N__29815),
            .in1(N__32247),
            .in2(N__30664),
            .in3(N__28485),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_20_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_20_4  (
            .in0(N__29819),
            .in1(N__32046),
            .in2(N__30677),
            .in3(N__27711),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_20_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_20_5  (
            .in0(N__29816),
            .in1(N__32607),
            .in2(N__30666),
            .in3(N__28272),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_20_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_20_6  (
            .in0(N__29818),
            .in1(N__32085),
            .in2(N__30676),
            .in3(N__27738),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_20_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_20_7  (
            .in0(N__29817),
            .in1(N__32411),
            .in2(N__30665),
            .in3(N__28122),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_21_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_21_0  (
            .in0(N__29803),
            .in1(N__32126),
            .in2(N__30688),
            .in3(N__28341),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_21_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_21_1  (
            .in0(N__29822),
            .in1(N__32373),
            .in2(N__30668),
            .in3(N__30834),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_3  (
            .in0(N__29823),
            .in1(N__32687),
            .in2(N__30670),
            .in3(N__27954),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_21_4 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_21_4  (
            .in0(N__32448),
            .in1(N__30588),
            .in2(N__29844),
            .in3(N__28086),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_21_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_10_21_5  (
            .in0(N__27837),
            .in1(N__29808),
            .in2(N__30669),
            .in3(N__32940),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_10_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_10_21_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_10_21_6  (
            .in0(N__29807),
            .in1(N__32939),
            .in2(N__30689),
            .in3(N__27836),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_22_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_22_3  (
            .in0(N__28212),
            .in1(N__29824),
            .in2(N__30671),
            .in3(N__32868),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_11_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_11_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_11_7_4 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \phase_controller_inst2.state_2_LC_11_7_4  (
            .in0(N__27439),
            .in1(N__31760),
            .in2(N__27472),
            .in3(N__40794),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46023),
            .ce(),
            .sr(N__45458));
    defparam \phase_controller_inst2.state_3_LC_11_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_11_8_1 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.state_3_LC_11_8_1  (
            .in0(N__27441),
            .in1(N__27504),
            .in2(N__27473),
            .in3(N__30969),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46015),
            .ce(),
            .sr(N__45465));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_11_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_11_9_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_9_LC_11_9_2  (
            .in0(N__33434),
            .in1(N__31996),
            .in2(_gnd_net_),
            .in3(N__31936),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_11_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_11_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__27462),
            .in2(_gnd_net_),
            .in3(N__27440),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_11_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_11_10_1 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_11_10_1  (
            .in0(N__33440),
            .in1(N__32001),
            .in2(_gnd_net_),
            .in3(N__31938),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45997),
            .ce(N__29320),
            .sr(N__45481));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_11_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_11_10_3 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_11_10_3  (
            .in0(N__28598),
            .in1(N__36368),
            .in2(N__31896),
            .in3(N__28687),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45997),
            .ce(N__29320),
            .sr(N__45481));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_11_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_11_10_4 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_11_10_4  (
            .in0(N__28686),
            .in1(N__31891),
            .in2(N__36488),
            .in3(N__28597),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45997),
            .ce(N__29320),
            .sr(N__45481));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_11_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_11_11_0 .LUT_INIT=16'b1010101011101111;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_11_11_0  (
            .in0(N__33384),
            .in1(N__31998),
            .in2(N__33132),
            .in3(N__31482),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_11_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_11_11_2 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_11_11_2  (
            .in0(N__35989),
            .in1(_gnd_net_),
            .in2(N__28691),
            .in3(N__31885),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_11_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_11_11_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_11_11_3  (
            .in0(N__31883),
            .in1(N__28671),
            .in2(_gnd_net_),
            .in3(N__35729),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_11_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_11_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__31480),
            .in2(_gnd_net_),
            .in3(N__33302),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_11_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_11_11_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_11_11_5  (
            .in0(N__31481),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33357),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_11_11_6 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_11_11_6  (
            .in0(N__28667),
            .in1(N__28619),
            .in2(N__35795),
            .in3(N__31884),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_11_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_11_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_11_11_7  (
            .in0(N__31997),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33433),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45986),
            .ce(N__29280),
            .sr(N__45486));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27653),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_12_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__29691),
            .in2(N__27531),
            .in3(N__29214),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32863),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32565),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_RNO_1_25_LC_11_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_RNO_1_25_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_RNO_1_25_LC_11_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_RNO_1_25_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__29690),
            .in2(_gnd_net_),
            .in3(N__30614),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29211),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_13_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_11_13_5  (
            .in0(N__29212),
            .in1(_gnd_net_),
            .in2(N__27663),
            .in3(N__30859),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32993),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45972),
            .ce(N__32965),
            .sr(N__45496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33695),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45972),
            .ce(N__32965),
            .sr(N__45496));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__27660),
            .in2(N__27654),
            .in3(N__27652),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__30735),
            .in2(_gnd_net_),
            .in3(N__27612),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__31689),
            .in2(_gnd_net_),
            .in3(N__27588),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__28716),
            .in2(_gnd_net_),
            .in3(N__27585),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__29433),
            .in2(_gnd_net_),
            .in3(N__27813),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__28710),
            .in2(_gnd_net_),
            .in3(N__27810),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__30741),
            .in2(_gnd_net_),
            .in3(N__27777),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__29415),
            .in2(_gnd_net_),
            .in3(N__27774),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__30789),
            .in2(_gnd_net_),
            .in3(N__27747),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__30795),
            .in2(_gnd_net_),
            .in3(N__27744),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__29427),
            .in2(_gnd_net_),
            .in3(N__27741),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__29421),
            .in2(_gnd_net_),
            .in3(N__27714),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__30765),
            .in2(_gnd_net_),
            .in3(N__27684),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__30777),
            .in2(_gnd_net_),
            .in3(N__27924),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__29409),
            .in2(_gnd_net_),
            .in3(N__27921),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__27918),
            .in2(_gnd_net_),
            .in3(N__27909),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__27906),
            .in2(_gnd_net_),
            .in3(N__27870),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__30981),
            .in2(_gnd_net_),
            .in3(N__27849),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__30993),
            .in2(_gnd_net_),
            .in3(N__27846),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__30783),
            .in2(_gnd_net_),
            .in3(N__27843),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_16_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31005),
            .in3(N__27840),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__30759),
            .in2(_gnd_net_),
            .in3(N__27816),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__30771),
            .in2(_gnd_net_),
            .in3(N__28014),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__28011),
            .in2(_gnd_net_),
            .in3(N__28002),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__30753),
            .in2(_gnd_net_),
            .in3(N__27984),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__30975),
            .in2(_gnd_net_),
            .in3(N__27981),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__30987),
            .in2(_gnd_net_),
            .in3(N__27960),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__30747),
            .in2(_gnd_net_),
            .in3(N__27957),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__28164),
            .in2(_gnd_net_),
            .in3(N__27930),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27927),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_11_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_11_17_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28227),
            .in3(N__29782),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_11_17_7  (
            .in0(N__29783),
            .in1(N__32856),
            .in2(N__30693),
            .in3(N__28205),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_18_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_11_18_0  (
            .in0(N__29813),
            .in1(N__28143),
            .in2(N__30605),
            .in3(N__32783),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_18_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_11_18_1  (
            .in0(N__32679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_18_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_11_18_3  (
            .in0(N__28142),
            .in1(N__29812),
            .in2(N__32784),
            .in3(N__30482),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_11_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_11_18_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_11_18_4  (
            .in0(N__29810),
            .in1(N__28141),
            .in2(_gnd_net_),
            .in3(N__32779),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_11_18_5  (
            .in0(N__29842),
            .in1(N__32412),
            .in2(N__30606),
            .in3(N__28118),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_11_18_6  (
            .in0(N__29811),
            .in1(N__32447),
            .in2(N__30604),
            .in3(N__28082),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_19_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_11_19_0  (
            .in0(N__29833),
            .in1(N__28046),
            .in2(N__30568),
            .in3(N__32907),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_11_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_11_19_2 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_11_19_2  (
            .in0(N__28481),
            .in1(N__30393),
            .in2(N__29846),
            .in3(N__32243),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_19_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_11_19_3  (
            .in0(N__30830),
            .in1(N__29832),
            .in2(N__30567),
            .in3(N__32369),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_19_4  (
            .in0(N__29828),
            .in1(N__31607),
            .in2(N__30569),
            .in3(N__28433),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_19_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_11_19_5  (
            .in0(N__29843),
            .in1(N__32724),
            .in2(N__30566),
            .in3(N__28404),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_20_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_11_20_1  (
            .in0(N__29836),
            .in1(N__32168),
            .in2(N__30686),
            .in3(N__28370),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_11_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_11_20_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_11_20_4  (
            .in0(N__30647),
            .in1(N__29837),
            .in2(N__32127),
            .in3(N__28337),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_20_5 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_11_20_5  (
            .in0(N__28304),
            .in1(N__30648),
            .in2(N__29847),
            .in3(N__32645),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_20_6 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_11_20_6  (
            .in0(N__28268),
            .in1(N__29841),
            .in2(N__30687),
            .in3(N__32606),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_11_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_11_21_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_11_21_0  (
            .in0(N__28584),
            .in1(N__29835),
            .in2(N__30691),
            .in3(N__32567),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_21_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_11_21_7  (
            .in0(N__29834),
            .in1(N__32566),
            .in2(N__30690),
            .in3(N__28583),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_11_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_11_22_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIF4PE_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__29845),
            .in2(_gnd_net_),
            .in3(N__28557),
            .lcout(\current_shift_inst.un4_control_input_0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__28501),
            .in2(_gnd_net_),
            .in3(N__37644),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_463_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_5_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_12_5_5  (
            .in0(N__33062),
            .in1(N__31077),
            .in2(N__45623),
            .in3(N__31094),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46033),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_12_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_6_3 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_12_6_3  (
            .in0(N__33068),
            .in1(N__31076),
            .in2(_gnd_net_),
            .in3(N__31093),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46022),
            .ce(),
            .sr(N__45452));
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_tr_sig_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_tr_sig_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33069),
            .lcout(\delay_measurement_inst.prev_tr_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46022),
            .ce(),
            .sr(N__45452));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_12_6_5 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_12_6_5  (
            .in0(N__28505),
            .in1(N__28518),
            .in2(_gnd_net_),
            .in3(N__37649),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46022),
            .ce(),
            .sr(N__45452));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_12_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_12_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__31759),
            .in2(_gnd_net_),
            .in3(N__40793),
            .lcout(\phase_controller_inst2.start_timer_hc_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_7_4 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_12_7_4  (
            .in0(N__28517),
            .in1(N__28506),
            .in2(_gnd_net_),
            .in3(N__37648),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_464_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_12_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_12_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_12_8_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_12_8_0  (
            .in0(N__28699),
            .in1(N__35948),
            .in2(_gnd_net_),
            .in3(N__31882),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46005),
            .ce(N__35369),
            .sr(N__45459));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_12_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_12_8_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_12_8_2  (
            .in0(N__28698),
            .in1(N__35997),
            .in2(_gnd_net_),
            .in3(N__31881),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46005),
            .ce(N__35369),
            .sr(N__45459));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_12_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43776),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46005),
            .ce(N__35369),
            .sr(N__45459));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_12_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_12_8_4 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_12_8_4  (
            .in0(N__28605),
            .in1(N__36372),
            .in2(N__28703),
            .in3(N__31880),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46005),
            .ce(N__35369),
            .sr(N__45459));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_12_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_12_8_5 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_12_8_5  (
            .in0(N__31879),
            .in1(N__28694),
            .in2(N__36489),
            .in3(N__28604),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46005),
            .ce(N__35369),
            .sr(N__45459));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_12_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_12_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_12_9_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_12_9_0  (
            .in0(N__32000),
            .in1(N__33435),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_12_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_12_9_1 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_12_9_1  (
            .in0(N__31875),
            .in1(N__28693),
            .in2(_gnd_net_),
            .in3(N__35733),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_12_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_12_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__31462),
            .in2(_gnd_net_),
            .in3(N__33303),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_12_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_12_9_3 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__31999),
            .in2(N__33441),
            .in3(N__31937),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_12_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_12_9_4 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_12_9_4  (
            .in0(N__28692),
            .in1(N__28623),
            .in2(N__35799),
            .in3(N__31877),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_12_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_12_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_12_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_12_9_5  (
            .in0(N__31876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35906),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_12_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_12_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__35840),
            .in2(_gnd_net_),
            .in3(N__31878),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_12_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_12_9_7  (
            .in0(N__31461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33257),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45996),
            .ce(N__35374),
            .sr(N__45466));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_12_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__31465),
            .in2(_gnd_net_),
            .in3(N__33356),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45985),
            .ce(N__35370),
            .sr(N__45473));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_12_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_12_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4_3_LC_12_11_0  (
            .in0(N__31917),
            .in1(N__35941),
            .in2(N__35996),
            .in3(N__31966),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_12_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0_6_LC_12_11_2  (
            .in0(N__28638),
            .in1(N__33127),
            .in2(_gnd_net_),
            .in3(N__31967),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a3_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_12_11_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1_6_LC_12_11_3  (
            .in0(N__35833),
            .in1(N__35899),
            .in2(_gnd_net_),
            .in3(N__35728),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_12_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_LC_12_11_4  (
            .in0(N__28632),
            .in1(N__33450),
            .in2(N__28626),
            .in3(N__33102),
            .lcout(\phase_controller_inst1.stoper_tr.N_257 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_12_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_12_11_5 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a3_1_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__36367),
            .in2(N__28608),
            .in3(N__35788),
            .lcout(\phase_controller_inst1.stoper_tr.N_240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_12_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a3_1_LC_12_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a3_1_LC_12_12_2  (
            .in0(N__29373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38217),
            .lcout(state_ns_i_a3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_12_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNIH19L_0_LC_12_12_3  (
            .in0(N__29104),
            .in1(N__28769),
            .in2(_gnd_net_),
            .in3(N__28887),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_13_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_13_3  (
            .in0(N__29581),
            .in1(N__31672),
            .in2(N__30674),
            .in3(N__29252),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_13_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_12_13_5  (
            .in0(N__29580),
            .in1(N__29220),
            .in2(_gnd_net_),
            .in3(N__29213),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_12_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_12_13_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_RNID9EC_0_LC_12_13_7  (
            .in0(N__28866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28751),
            .lcout(\phase_controller_inst2.stoper_tr.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_14_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_0_LC_12_14_0  (
            .in0(N__28767),
            .in1(N__28883),
            .in2(N__29115),
            .in3(N__29159),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45962),
            .ce(N__42507),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_14_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.stoper_state_1_LC_12_14_1  (
            .in0(N__29160),
            .in1(N__29111),
            .in2(N__28927),
            .in3(N__28768),
            .lcout(\phase_controller_inst2.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45962),
            .ce(N__42507),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31590),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32313),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_12_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_12_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32268),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31657),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_12_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_12_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_12_15_1  (
            .in0(N__29799),
            .in1(N__31550),
            .in2(N__30675),
            .in3(N__30722),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_15_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_12_15_2  (
            .in0(N__30615),
            .in1(N__29800),
            .in2(N__32336),
            .in3(N__29466),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31549),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32101),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_12_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32067),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_12_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32227),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_12_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_12_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32587),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32148),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32187),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32394),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32626),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32889),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32022),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_12_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32923),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32803),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32707),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32356),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32428),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32740),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32464),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32771),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_12_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_18_6 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_18_6  (
            .in0(N__30968),
            .in1(N__36149),
            .in2(N__36115),
            .in3(N__37623),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45947),
            .ce(),
            .sr(N__45531));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_12_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_12_18_7  (
            .in0(N__30948),
            .in1(N__32357),
            .in2(_gnd_net_),
            .in3(N__30829),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_19_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_19_0  (
            .in0(N__31159),
            .in1(N__31187),
            .in2(_gnd_net_),
            .in3(N__31137),
            .lcout(\current_shift_inst.timer_s1.N_186_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31158),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__36095),
            .in2(_gnd_net_),
            .in3(N__36148),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_LC_12_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_12_20_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_12_20_2  (
            .in0(N__31186),
            .in1(N__31160),
            .in2(_gnd_net_),
            .in3(N__31136),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45940),
            .ce(),
            .sr(N__45543));
    defparam \current_shift_inst.start_timer_s1_LC_12_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_12_21_1 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_12_21_1  (
            .in0(N__33007),
            .in1(N__31182),
            .in2(_gnd_net_),
            .in3(N__36110),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45937),
            .ce(),
            .sr(N__45552));
    defparam \current_shift_inst.stop_timer_s1_LC_12_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_12_21_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_12_21_4  (
            .in0(N__36111),
            .in1(N__33008),
            .in2(N__31188),
            .in3(N__31135),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45937),
            .ce(),
            .sr(N__45552));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_12_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_12_22_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_12_22_1  (
            .in0(N__31161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31131),
            .lcout(\current_shift_inst.timer_s1.N_185_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.tr_state_0_LC_13_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.tr_state_0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.tr_state_0_LC_13_6_0 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \delay_measurement_inst.tr_state_0_LC_13_6_0  (
            .in0(N__33061),
            .in1(N__31075),
            .in2(_gnd_net_),
            .in3(N__31095),
            .lcout(\delay_measurement_inst.tr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46034),
            .ce(N__42508),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_13_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_13_7_0 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_13_7_0  (
            .in0(N__31059),
            .in1(N__38231),
            .in2(N__44559),
            .in3(N__31044),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46024),
            .ce(),
            .sr(N__45453));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1_c_inv_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__31038),
            .in2(N__31032),
            .in3(N__35311),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2_c_inv_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__31011),
            .in2(N__31023),
            .in3(N__35294),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3_c_inv_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__31305),
            .in2(N__31314),
            .in3(N__35261),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4_c_inv_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__31287),
            .in2(N__31299),
            .in3(N__35237),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5_c_inv_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__31272),
            .in2(N__31281),
            .in3(N__35510),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6_c_inv_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__31257),
            .in2(N__31266),
            .in3(N__35486),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7_c_inv_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__31239),
            .in2(N__31251),
            .in3(N__42197),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8_c_inv_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__31218),
            .in2(N__31233),
            .in3(N__42155),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9_c_inv_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__31212),
            .in2(N__31506),
            .in3(N__42119),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_9_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10_c_inv_LC_13_9_1  (
            .in0(N__35456),
            .in1(N__31194),
            .in2(N__31206),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11_c_inv_LC_13_9_2  (
            .in0(N__35435),
            .in1(N__31416),
            .in2(N__31428),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12_c_inv_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__31398),
            .in2(N__31410),
            .in3(N__35414),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13_c_inv_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__31383),
            .in2(N__31392),
            .in3(N__35654),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14_c_inv_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__31365),
            .in2(N__31377),
            .in3(N__35630),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15_c_inv_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__31350),
            .in2(N__31359),
            .in3(N__35609),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16_c_inv_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__31344),
            .in2(N__31494),
            .in3(N__38118),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17_c_inv_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__31326),
            .in2(N__31338),
            .in3(N__35579),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_17 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18_c_inv_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__31320),
            .in2(N__31524),
            .in3(N__35555),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_inv_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__31533),
            .in2(N__31515),
            .in3(N__35534),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31527),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43556),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45998),
            .ce(N__35379),
            .sr(N__45467));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38037),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45998),
            .ce(N__35379),
            .sr(N__45467));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_13_11_4 .LUT_INIT=16'b1111111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_13_11_4  (
            .in0(N__31478),
            .in1(N__31979),
            .in2(N__33131),
            .in3(N__33377),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45987),
            .ce(N__35378),
            .sr(N__45474));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_13_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_13_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38075),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45987),
            .ce(N__35378),
            .sr(N__45474));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_11_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__31479),
            .in2(_gnd_net_),
            .in3(N__33320),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45987),
            .ce(N__35378),
            .sr(N__45474));
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_13_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_14_LC_13_12_0 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_14_LC_13_12_0  (
            .in0(N__38511),
            .in1(N__43661),
            .in2(N__31809),
            .in3(N__43728),
            .lcout(measured_delay_tr_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45978),
            .ce(N__43520),
            .sr(N__45482));
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_12_1 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_15_LC_13_12_1  (
            .in0(N__43729),
            .in1(N__37994),
            .in2(N__43676),
            .in3(N__38460),
            .lcout(measured_delay_tr_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45978),
            .ce(N__43520),
            .sr(N__45482));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_12_6 .LUT_INIT=16'b1111010111110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2_6_LC_13_12_6  (
            .in0(N__31971),
            .in1(N__31918),
            .in2(N__33439),
            .in3(N__33101),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_o2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_13_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_13_12_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_14_LC_13_12_7  (
            .in0(N__43660),
            .in1(N__37993),
            .in2(_gnd_net_),
            .in3(N__38459),
            .lcout(\delay_measurement_inst.delay_tr_reg_esr_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_13_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNITN7V_0_LC_13_13_2  (
            .in0(N__43285),
            .in1(N__43083),
            .in2(_gnd_net_),
            .in3(N__43429),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_1_LC_13_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_13_14_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_1_LC_13_14_0  (
            .in0(N__31800),
            .in1(N__31770),
            .in2(N__31726),
            .in3(N__40792),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45968),
            .ce(),
            .sr(N__45490));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31624),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__33696),
            .in2(N__33632),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__33605),
            .in2(N__33665),
            .in3(N__31611),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__33584),
            .in2(N__33633),
            .in3(N__31569),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__33606),
            .in2(N__33563),
            .in3(N__31536),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__33585),
            .in2(N__33537),
            .in3(N__32295),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__33503),
            .in2(N__33564),
            .in3(N__32250),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__33533),
            .in2(N__33476),
            .in3(N__32211),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__33504),
            .in2(N__33902),
            .in3(N__32172),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__45963),
            .ce(N__32964),
            .sr(N__45497));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__33872),
            .in2(N__33480),
            .in3(N__32130),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__33845),
            .in2(N__33909),
            .in3(N__32088),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__33824),
            .in2(N__33876),
            .in3(N__32049),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__33846),
            .in2(N__33803),
            .in3(N__32004),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__33825),
            .in2(N__33776),
            .in3(N__32610),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__33746),
            .in2(N__33804),
            .in3(N__32571),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__33715),
            .in2(N__33777),
            .in3(N__32529),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__33747),
            .in2(N__34145),
            .in3(N__32487),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__45957),
            .ce(N__32963),
            .sr(N__45506));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__34118),
            .in2(N__33723),
            .in3(N__32451),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__34094),
            .in2(N__34152),
            .in3(N__32415),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__34119),
            .in2(N__34073),
            .in3(N__32376),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__34095),
            .in2(N__34043),
            .in3(N__32340),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__34016),
            .in2(N__34074),
            .in3(N__32910),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__33995),
            .in2(N__34044),
            .in3(N__32871),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__34017),
            .in2(N__33962),
            .in3(N__32826),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__33925),
            .in2(N__33996),
            .in3(N__32787),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__45953),
            .ce(N__32962),
            .sr(N__45514));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__34922),
            .in2(N__33966),
            .in3(N__32760),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__45950),
            .ce(N__32961),
            .sr(N__45523));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__34895),
            .in2(N__33936),
            .in3(N__32727),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__45950),
            .ce(N__32961),
            .sr(N__45523));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__34875),
            .in2(N__34926),
            .in3(N__32691),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__45950),
            .ce(N__32961),
            .sr(N__45523));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__34896),
            .in2(N__34719),
            .in3(N__32652),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__45950),
            .ce(N__32961),
            .sr(N__45523));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32649),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32978),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45950),
            .ce(N__32961),
            .sr(N__45523));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_19_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_13_19_1  (
            .in0(N__43114),
            .in1(N__43470),
            .in2(N__43338),
            .in3(N__36504),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45948),
            .ce(),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_19_3 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_13_19_3  (
            .in0(N__43115),
            .in1(N__43471),
            .in2(N__43339),
            .in3(N__36294),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45948),
            .ce(),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_19_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_13_19_4  (
            .in0(N__43468),
            .in1(N__43316),
            .in2(N__43127),
            .in3(N__36246),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45948),
            .ce(),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_19_5 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_13_19_5  (
            .in0(N__43116),
            .in1(N__36213),
            .in2(N__43340),
            .in3(N__43473),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45948),
            .ce(),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_19_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_13_19_6  (
            .in0(N__43469),
            .in1(N__43317),
            .in2(N__43128),
            .in3(N__36180),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45948),
            .ce(),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_19_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_13_19_7  (
            .in0(N__43117),
            .in1(N__43472),
            .in2(N__43341),
            .in3(N__36618),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45948),
            .ce(),
            .sr(N__45532));
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_13_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_0_LC_13_20_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_0_LC_13_20_0  (
            .in0(N__42078),
            .in1(N__41522),
            .in2(N__46941),
            .in3(N__41750),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_13_20_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_13_20_1  (
            .in0(N__41747),
            .in1(N__46918),
            .in2(N__41538),
            .in3(N__40991),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_13_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_13_20_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_13_20_2  (
            .in0(N__41123),
            .in1(N__41525),
            .in2(N__46944),
            .in3(N__41753),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_13_20_3 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_13_20_3  (
            .in0(N__41521),
            .in1(N__46754),
            .in2(N__41376),
            .in3(N__46921),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_13_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_13_20_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_13_20_4  (
            .in0(N__41071),
            .in1(N__41523),
            .in2(N__46942),
            .in3(N__41751),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_13_20_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_13_20_5  (
            .in0(N__41749),
            .in1(N__46920),
            .in2(N__41540),
            .in3(N__40945),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_13_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_13_20_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_13_20_6  (
            .in0(N__41034),
            .in1(N__41524),
            .in2(N__46943),
            .in3(N__41752),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_13_20_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_13_20_7  (
            .in0(N__41748),
            .in1(N__46919),
            .in2(N__41539),
            .in3(N__41816),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45945),
            .ce(N__38932),
            .sr(N__45539));
    defparam \phase_controller_inst1.S1_LC_13_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36116),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45941),
            .ce(),
            .sr(N__45544));
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_13_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_13_22_1 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_3_LC_13_22_1 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_3_LC_13_22_1  (
            .in0(N__46274),
            .in1(N__42401),
            .in2(N__46498),
            .in3(N__41622),
            .lcout(measured_delay_hc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45938),
            .ce(),
            .sr(N__45553));
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_13_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_8_LC_13_22_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_8_LC_13_22_2  (
            .in0(N__39530),
            .in1(N__46481),
            .in2(N__40937),
            .in3(N__46275),
            .lcout(measured_delay_hc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45938),
            .ce(),
            .sr(N__45553));
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_13_LC_13_22_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_13_LC_13_22_4  (
            .in0(N__39240),
            .in1(N__46473),
            .in2(N__41817),
            .in3(N__46271),
            .lcout(measured_delay_hc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45938),
            .ce(),
            .sr(N__45553));
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_13_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_13_22_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_21_LC_13_22_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_21_LC_13_22_6  (
            .in0(N__39554),
            .in1(N__46474),
            .in2(_gnd_net_),
            .in3(N__46272),
            .lcout(measured_delay_hc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45938),
            .ce(),
            .sr(N__45553));
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_22_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_22_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_22_LC_13_22_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_22_LC_13_22_7  (
            .in0(N__46273),
            .in1(_gnd_net_),
            .in2(N__46497),
            .in3(N__39173),
            .lcout(measured_delay_hc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45938),
            .ce(),
            .sr(N__45553));
    defparam SB_DFF_inst_DELAY_TR1_LC_14_5_0.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR1_LC_14_5_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR1_LC_14_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR1_LC_14_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33087),
            .lcout(delay_tr_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46051),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_TR2_LC_14_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_TR2_LC_14_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_TR2_LC_14_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_TR2_LC_14_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33075),
            .lcout(delay_tr_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46051),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_14_5_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_14_5_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_14_5_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_14_5_6 (
            .in0(N__33042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46051),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_7_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_0_LC_14_7_3  (
            .in0(N__42630),
            .in1(N__42797),
            .in2(N__42960),
            .in3(N__42673),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46035),
            .ce(N__42509),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_8_0 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_8_0  (
            .in0(N__42621),
            .in1(N__42951),
            .in2(N__42805),
            .in3(N__35445),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_8_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_1_LC_14_8_1  (
            .in0(N__38156),
            .in1(N__35315),
            .in2(_gnd_net_),
            .in3(N__42672),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_8_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_8_2  (
            .in0(N__42624),
            .in1(N__42950),
            .in2(N__33024),
            .in3(N__42780),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_8_3 .LUT_INIT=16'b1010100010100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_8_3  (
            .in0(N__35424),
            .in1(N__42625),
            .in2(N__42808),
            .in3(N__42947),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_8_4 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_8_4  (
            .in0(N__42622),
            .in1(N__42952),
            .in2(N__42806),
            .in3(N__35403),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_8_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_8_5  (
            .in0(N__42948),
            .in1(N__42626),
            .in2(N__35643),
            .in3(N__42775),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_8_6 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_8_6  (
            .in0(N__42623),
            .in1(N__42953),
            .in2(N__42807),
            .in3(N__35619),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_8_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_8_7  (
            .in0(N__42949),
            .in1(N__42627),
            .in2(N__35598),
            .in3(N__42776),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46025),
            .ce(),
            .sr(N__45454));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_9_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_9_0  (
            .in0(N__42603),
            .in1(N__42934),
            .in2(N__35568),
            .in3(N__42789),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_9_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_9_1  (
            .in0(N__42785),
            .in1(N__42607),
            .in2(N__42955),
            .in3(N__35544),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_9_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_9_2  (
            .in0(N__42604),
            .in1(N__42935),
            .in2(N__35520),
            .in3(N__42790),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_9_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_9_3  (
            .in0(N__42786),
            .in1(N__42608),
            .in2(N__42956),
            .in3(N__35283),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_9_4 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_9_4  (
            .in0(N__42605),
            .in1(N__42936),
            .in2(N__35250),
            .in3(N__42791),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_9_5 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_9_5  (
            .in0(N__42787),
            .in1(N__42609),
            .in2(N__42957),
            .in3(N__35226),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_9_6 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_9_6  (
            .in0(N__42606),
            .in1(N__42937),
            .in2(N__35499),
            .in3(N__42792),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_9_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_9_7  (
            .in0(N__42788),
            .in1(N__42610),
            .in2(N__42958),
            .in3(N__35475),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46016),
            .ce(),
            .sr(N__45456));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_14_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_14_10_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_14_10_2  (
            .in0(N__33231),
            .in1(N__33204),
            .in2(_gnd_net_),
            .in3(N__33177),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOE_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(N__38149),
            .in2(_gnd_net_),
            .in3(N__42659),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19_c_RNICDOEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_14_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_14_10_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIBL28_0_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(N__42581),
            .in2(_gnd_net_),
            .in3(N__42781),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed11 ),
            .ltout(\phase_controller_inst1.stoper_tr.time_passed11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33135),
            .in3(N__42658),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_15_LC_14_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_15_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_15_LC_14_11_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_15_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__45618),
            .in2(_gnd_net_),
            .in3(N__36415),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_14_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_14_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0_6_LC_14_11_2  (
            .in0(N__33289),
            .in1(N__33319),
            .in2(N__33250),
            .in3(N__33343),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_14_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_14_11_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2_9_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33105),
            .in3(N__33376),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f1_0_i_i_a2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_14_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_14_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3_3_LC_14_11_5  (
            .in0(N__43542),
            .in1(N__43761),
            .in2(N__38041),
            .in3(N__38073),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_f0_0_a2_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_14_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_14_11_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_i_o2_15_LC_14_11_7  (
            .in0(N__43543),
            .in1(N__43762),
            .in2(N__38042),
            .in3(N__38074),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_6_i_o2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_14_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_14_12_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_RNO_0_9_LC_14_12_0  (
            .in0(N__38627),
            .in1(N__43707),
            .in2(N__38469),
            .in3(N__35685),
            .lcout(),
            .ltout(\delay_measurement_inst.N_360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_14_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_9_LC_14_12_1 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_9_LC_14_12_1  (
            .in0(N__38628),
            .in1(N__33273),
            .in2(N__33387),
            .in3(N__43671),
            .lcout(measured_delay_tr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45988),
            .ce(N__43519),
            .sr(N__45475));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_14_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_14_12_2 .LUT_INIT=16'b1111111100001110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM4EJ7_14_LC_14_12_2  (
            .in0(N__38464),
            .in1(N__38510),
            .in2(N__37995),
            .in3(N__43706),
            .lcout(\delay_measurement_inst.N_354 ),
            .ltout(\delay_measurement_inst.N_354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_14_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_10_LC_14_12_3 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_10_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(N__43665),
            .in2(N__33360),
            .in3(N__38589),
            .lcout(measured_delay_tr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45988),
            .ce(N__43519),
            .sr(N__45475));
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_14_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_11_LC_14_12_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_11_LC_14_12_5  (
            .in0(N__38568),
            .in1(N__43666),
            .in2(_gnd_net_),
            .in3(N__33270),
            .lcout(measured_delay_tr_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45988),
            .ce(N__43519),
            .sr(N__45475));
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_14_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_12_LC_14_12_6 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_12_LC_14_12_6  (
            .in0(N__33271),
            .in1(_gnd_net_),
            .in2(N__43677),
            .in3(N__38550),
            .lcout(measured_delay_tr_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45988),
            .ce(N__43519),
            .sr(N__45475));
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_14_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_14_12_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_13_LC_14_12_7 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_13_LC_14_12_7  (
            .in0(N__38532),
            .in1(N__33272),
            .in2(_gnd_net_),
            .in3(N__43670),
            .lcout(measured_delay_tr_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45988),
            .ce(N__43519),
            .sr(N__45475));
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_14_13_0  (
            .in0(N__34842),
            .in1(N__33688),
            .in2(_gnd_net_),
            .in3(N__33669),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_14_13_1  (
            .in0(N__34850),
            .in1(N__33652),
            .in2(_gnd_net_),
            .in3(N__33636),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_14_13_2  (
            .in0(N__34843),
            .in1(N__33625),
            .in2(_gnd_net_),
            .in3(N__33609),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_14_13_3  (
            .in0(N__34851),
            .in1(N__33604),
            .in2(_gnd_net_),
            .in3(N__33588),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_14_13_4  (
            .in0(N__34844),
            .in1(N__33583),
            .in2(_gnd_net_),
            .in3(N__33567),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_14_13_5  (
            .in0(N__34852),
            .in1(N__33556),
            .in2(_gnd_net_),
            .in3(N__33540),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_14_13_6  (
            .in0(N__34845),
            .in1(N__33529),
            .in2(_gnd_net_),
            .in3(N__33507),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_14_13_7  (
            .in0(N__34853),
            .in1(N__33497),
            .in2(_gnd_net_),
            .in3(N__33483),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__45979),
            .ce(N__34700),
            .sr(N__45483));
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_14_14_0  (
            .in0(N__34841),
            .in1(N__33475),
            .in2(_gnd_net_),
            .in3(N__33453),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_14_14_1  (
            .in0(N__34837),
            .in1(N__33901),
            .in2(_gnd_net_),
            .in3(N__33879),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_14_14_2  (
            .in0(N__34838),
            .in1(N__33865),
            .in2(_gnd_net_),
            .in3(N__33849),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_14_14_3  (
            .in0(N__34834),
            .in1(N__33844),
            .in2(_gnd_net_),
            .in3(N__33828),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_14_14_4  (
            .in0(N__34839),
            .in1(N__33823),
            .in2(_gnd_net_),
            .in3(N__33807),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_14_14_5  (
            .in0(N__34835),
            .in1(N__33796),
            .in2(_gnd_net_),
            .in3(N__33780),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_14_14_6  (
            .in0(N__34840),
            .in1(N__33764),
            .in2(_gnd_net_),
            .in3(N__33750),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_14_14_7  (
            .in0(N__34836),
            .in1(N__33740),
            .in2(_gnd_net_),
            .in3(N__33726),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__45973),
            .ce(N__34701),
            .sr(N__45487));
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_14_15_0  (
            .in0(N__34846),
            .in1(N__33719),
            .in2(_gnd_net_),
            .in3(N__33699),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_14_15_1  (
            .in0(N__34854),
            .in1(N__34144),
            .in2(_gnd_net_),
            .in3(N__34122),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_14_15_2  (
            .in0(N__34847),
            .in1(N__34112),
            .in2(_gnd_net_),
            .in3(N__34098),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_14_15_3  (
            .in0(N__34855),
            .in1(N__34093),
            .in2(_gnd_net_),
            .in3(N__34077),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_14_15_4  (
            .in0(N__34848),
            .in1(N__34061),
            .in2(_gnd_net_),
            .in3(N__34047),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_14_15_5  (
            .in0(N__34856),
            .in1(N__34036),
            .in2(_gnd_net_),
            .in3(N__34020),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_14_15_6  (
            .in0(N__34849),
            .in1(N__34015),
            .in2(_gnd_net_),
            .in3(N__33999),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_14_15_7  (
            .in0(N__34857),
            .in1(N__33988),
            .in2(_gnd_net_),
            .in3(N__33969),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__45969),
            .ce(N__34696),
            .sr(N__45491));
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_14_16_0  (
            .in0(N__34830),
            .in1(N__33961),
            .in2(_gnd_net_),
            .in3(N__33939),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__45964),
            .ce(N__34695),
            .sr(N__45498));
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_14_16_1  (
            .in0(N__34774),
            .in1(N__33929),
            .in2(_gnd_net_),
            .in3(N__34929),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__45964),
            .ce(N__34695),
            .sr(N__45498));
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_14_16_2  (
            .in0(N__34831),
            .in1(N__34915),
            .in2(_gnd_net_),
            .in3(N__34899),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__45964),
            .ce(N__34695),
            .sr(N__45498));
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_14_16_3  (
            .in0(N__34775),
            .in1(N__34894),
            .in2(_gnd_net_),
            .in3(N__34878),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__45964),
            .ce(N__34695),
            .sr(N__45498));
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_14_16_4  (
            .in0(N__34832),
            .in1(N__34874),
            .in2(_gnd_net_),
            .in3(N__34860),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__45964),
            .ce(N__34695),
            .sr(N__45498));
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_16_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_14_16_5  (
            .in0(N__34715),
            .in1(N__34833),
            .in2(_gnd_net_),
            .in3(N__34722),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45964),
            .ce(N__34695),
            .sr(N__45498));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_14_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_14_17_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_14_17_0  (
            .in0(N__41940),
            .in1(N__40902),
            .in2(N__41541),
            .in3(N__46934),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45958),
            .ce(N__38925),
            .sr(N__45507));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_17_6  (
            .in0(N__34653),
            .in1(N__34574),
            .in2(_gnd_net_),
            .in3(N__34629),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_17_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_17_7  (
            .in0(N__34575),
            .in1(_gnd_net_),
            .in2(N__34209),
            .in3(N__34205),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_18_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_18_0  (
            .in0(N__43098),
            .in1(N__43446),
            .in2(N__43331),
            .in3(N__36579),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45954),
            .ce(),
            .sr(N__45515));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_14_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_14_18_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_1_LC_14_18_1  (
            .in0(N__43156),
            .in1(N__39098),
            .in2(_gnd_net_),
            .in3(N__36332),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_14_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_14_18_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_14_18_2  (
            .in0(N__43290),
            .in1(N__43101),
            .in2(N__34962),
            .in3(N__43449),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45954),
            .ce(),
            .sr(N__45515));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_18_3 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_18_3  (
            .in0(N__43444),
            .in1(N__43291),
            .in2(N__43124),
            .in3(N__36555),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45954),
            .ce(),
            .sr(N__45515));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_18_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_18_4  (
            .in0(N__43099),
            .in1(N__43447),
            .in2(N__43332),
            .in3(N__36531),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45954),
            .ce(),
            .sr(N__45515));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_18_6 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_18_6  (
            .in0(N__43100),
            .in1(N__43448),
            .in2(N__43333),
            .in3(N__36735),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45954),
            .ce(),
            .sr(N__45515));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_18_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_18_7  (
            .in0(N__43445),
            .in1(N__43292),
            .in2(N__43125),
            .in3(N__36711),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45954),
            .ce(),
            .sr(N__45515));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_14_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_14_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__34959),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_14_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_14_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__34941),
            .in2(N__34953),
            .in3(N__36328),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_14_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_14_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__34935),
            .in2(N__39039),
            .in3(N__36305),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_14_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_14_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__35046),
            .in2(N__38952),
            .in3(N__36272),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_14_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_14_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__35031),
            .in2(N__35040),
            .in3(N__36224),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_14_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_14_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__35025),
            .in2(N__38979),
            .in3(N__36191),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_14_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_14_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__35019),
            .in2(N__38967),
            .in3(N__36629),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_14_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_14_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__35013),
            .in2(N__39027),
            .in3(N__38871),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_14_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_14_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__35007),
            .in2(N__35001),
            .in3(N__38847),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_14_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_14_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__34983),
            .in2(N__34992),
            .in3(N__36860),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_14_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_14_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__34968),
            .in2(N__34977),
            .in3(N__36594),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_14_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_14_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__35112),
            .in2(N__35124),
            .in3(N__36570),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_14_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_14_20_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_14_20_4  (
            .in0(N__36546),
            .in1(N__35097),
            .in2(N__35106),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_14_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_14_20_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_14_20_5  (
            .in0(N__36515),
            .in1(N__35082),
            .in2(N__35091),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_14_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_14_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__35076),
            .in2(N__38994),
            .in3(N__36750),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_14_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_14_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__35070),
            .in2(N__39012),
            .in3(N__36726),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_14_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_14_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__35064),
            .in2(N__36822),
            .in3(N__36702),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_14_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_14_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__35058),
            .in2(N__36813),
            .in3(N__36884),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_14_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_14_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__35052),
            .in2(N__36804),
            .in3(N__36842),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_14_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_14_21_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_14_21_3  (
            .in0(N__36647),
            .in1(N__35136),
            .in2(N__36831),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35130),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_14_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_14_21_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9K_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35127),
            .in3(N__39097),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19_c_RNIRS9KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_14_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_9_LC_14_22_2 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_9_LC_14_22_2  (
            .in0(N__46270),
            .in1(N__41360),
            .in2(N__46496),
            .in3(N__39138),
            .lcout(measured_delay_hc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45942),
            .ce(),
            .sr(N__45545));
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_14_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_14_LC_14_22_3 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_14_LC_14_22_3  (
            .in0(N__39156),
            .in1(N__46465),
            .in2(N__41592),
            .in3(N__46267),
            .lcout(measured_delay_hc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45942),
            .ce(),
            .sr(N__45545));
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_14_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_14_22_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_23_LC_14_22_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_23_LC_14_22_4  (
            .in0(N__46268),
            .in1(_gnd_net_),
            .in2(N__46495),
            .in3(N__39188),
            .lcout(measured_delay_hc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45942),
            .ce(),
            .sr(N__45545));
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_14_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_14_22_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_24_LC_14_22_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_24_LC_14_22_5  (
            .in0(N__39203),
            .in1(N__46469),
            .in2(_gnd_net_),
            .in3(N__46269),
            .lcout(measured_delay_hc_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45942),
            .ce(),
            .sr(N__45545));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBOIH1_14_LC_14_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBOIH1_14_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBOIH1_14_LC_14_23_1 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBOIH1_14_LC_14_23_1  (
            .in0(N__46292),
            .in1(N__39154),
            .in2(N__42400),
            .in3(N__39136),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_24_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_14_24_1  (
            .in0(_gnd_net_),
            .in1(N__36794),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45934),
            .ce(N__37856),
            .sr(N__45558));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_14_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_14_24_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_14_24_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_14_24_6  (
            .in0(_gnd_net_),
            .in1(N__36773),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45934),
            .ce(N__37856),
            .sr(N__45558));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_25_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_14_25_0  (
            .in0(N__37772),
            .in1(N__36790),
            .in2(_gnd_net_),
            .in3(N__35163),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_25_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_25_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_25_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_14_25_1  (
            .in0(N__37768),
            .in1(N__36769),
            .in2(_gnd_net_),
            .in3(N__35160),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_25_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_14_25_2  (
            .in0(N__37773),
            .in1(N__37111),
            .in2(_gnd_net_),
            .in3(N__35157),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_25_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_25_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_14_25_3  (
            .in0(N__37769),
            .in1(N__37079),
            .in2(_gnd_net_),
            .in3(N__35154),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_25_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_25_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_14_25_4  (
            .in0(N__37774),
            .in1(N__37055),
            .in2(_gnd_net_),
            .in3(N__35151),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_25_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_25_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_14_25_5  (
            .in0(N__37770),
            .in1(N__37031),
            .in2(_gnd_net_),
            .in3(N__35148),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_25_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_25_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_14_25_6  (
            .in0(N__37775),
            .in1(N__37001),
            .in2(_gnd_net_),
            .in3(N__35145),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_25_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_25_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_14_25_7  (
            .in0(N__37771),
            .in1(N__36971),
            .in2(_gnd_net_),
            .in3(N__35142),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__45933),
            .ce(N__37818),
            .sr(N__45564));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_26_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_26_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_14_26_0  (
            .in0(N__37736),
            .in1(N__36943),
            .in2(_gnd_net_),
            .in3(N__35139),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_26_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_26_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_26_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_14_26_1  (
            .in0(N__37726),
            .in1(N__36913),
            .in2(_gnd_net_),
            .in3(N__35190),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_26_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_26_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_14_26_2  (
            .in0(N__37733),
            .in1(N__37357),
            .in2(_gnd_net_),
            .in3(N__35187),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_26_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_26_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_14_26_3  (
            .in0(N__37723),
            .in1(N__37325),
            .in2(_gnd_net_),
            .in3(N__35184),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_26_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_26_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_14_26_4  (
            .in0(N__37734),
            .in1(N__37306),
            .in2(_gnd_net_),
            .in3(N__35181),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_26_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_14_26_5  (
            .in0(N__37724),
            .in1(N__37280),
            .in2(_gnd_net_),
            .in3(N__35178),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_26_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_26_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_14_26_6  (
            .in0(N__37735),
            .in1(N__37250),
            .in2(_gnd_net_),
            .in3(N__35175),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_26_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_26_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_26_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_14_26_7  (
            .in0(N__37725),
            .in1(N__37220),
            .in2(_gnd_net_),
            .in3(N__35172),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__45931),
            .ce(N__37810),
            .sr(N__45568));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_27_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_27_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_14_27_0  (
            .in0(N__37776),
            .in1(N__37195),
            .in2(_gnd_net_),
            .in3(N__35169),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_27_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_27_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_27_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_14_27_1  (
            .in0(N__37764),
            .in1(N__37165),
            .in2(_gnd_net_),
            .in3(N__35166),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_27_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_27_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_14_27_2  (
            .in0(N__37777),
            .in1(N__37135),
            .in2(_gnd_net_),
            .in3(N__35217),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_27_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_27_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_14_27_3  (
            .in0(N__37765),
            .in1(N__37595),
            .in2(_gnd_net_),
            .in3(N__35214),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_27_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_27_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_14_27_4  (
            .in0(N__37778),
            .in1(N__37571),
            .in2(_gnd_net_),
            .in3(N__35211),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_27_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_27_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_27_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_14_27_5  (
            .in0(N__37766),
            .in1(N__37547),
            .in2(_gnd_net_),
            .in3(N__35208),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_27_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_27_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_27_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_14_27_6  (
            .in0(N__37779),
            .in1(N__37517),
            .in2(_gnd_net_),
            .in3(N__35205),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_27_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_27_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_27_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_14_27_7  (
            .in0(N__37767),
            .in1(N__37487),
            .in2(_gnd_net_),
            .in3(N__35202),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__45929),
            .ce(N__37811),
            .sr(N__45571));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_28_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_28_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_28_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_14_28_0  (
            .in0(N__37727),
            .in1(N__37462),
            .in2(_gnd_net_),
            .in3(N__35199),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__45928),
            .ce(N__37809),
            .sr(N__45574));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_28_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_28_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_28_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_14_28_1  (
            .in0(N__37731),
            .in1(N__37432),
            .in2(_gnd_net_),
            .in3(N__35196),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__45928),
            .ce(N__37809),
            .sr(N__45574));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_28_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_28_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_28_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_14_28_2  (
            .in0(N__37728),
            .in1(N__37384),
            .in2(_gnd_net_),
            .in3(N__35193),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__45928),
            .ce(N__37809),
            .sr(N__45574));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_28_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_28_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_28_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_14_28_3  (
            .in0(N__37732),
            .in1(N__37882),
            .in2(_gnd_net_),
            .in3(N__35394),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__45928),
            .ce(N__37809),
            .sr(N__45574));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_28_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_28_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_28_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_14_28_4  (
            .in0(N__37729),
            .in1(N__37406),
            .in2(_gnd_net_),
            .in3(N__35391),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__45928),
            .ce(N__37809),
            .sr(N__45574));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_28_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_28_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_28_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_14_28_5  (
            .in0(N__37904),
            .in1(N__37730),
            .in2(_gnd_net_),
            .in3(N__35388),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45928),
            .ce(N__37809),
            .sr(N__45574));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_15_6_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_15_6_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_15_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_15_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35385),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46052),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_15_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_15_7_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_RNIEUJM_0_LC_15_7_5  (
            .in0(N__42848),
            .in1(N__42620),
            .in2(_gnd_net_),
            .in3(N__42753),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0_0_c_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__35325),
            .in2(N__35316),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_15_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_15_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_2_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__35295),
            .in2(_gnd_net_),
            .in3(N__35277),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_15_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_15_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_3_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__35274),
            .in2(N__35265),
            .in3(N__35241),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_15_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_15_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_4_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__35238),
            .in2(_gnd_net_),
            .in3(N__35220),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_15_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_15_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_5_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__35511),
            .in2(_gnd_net_),
            .in3(N__35490),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_15_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_15_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_6_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__35487),
            .in2(_gnd_net_),
            .in3(N__35469),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_15_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_15_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_7_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__42198),
            .in2(_gnd_net_),
            .in3(N__35466),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_15_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_15_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_8_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__42156),
            .in2(_gnd_net_),
            .in3(N__35463),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_15_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_15_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_9_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__42120),
            .in2(_gnd_net_),
            .in3(N__35460),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_9 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_15_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_15_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_10_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__35457),
            .in2(_gnd_net_),
            .in3(N__35439),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_15_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_15_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_11_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__35436),
            .in2(_gnd_net_),
            .in3(N__35418),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_15_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_15_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_12_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__35415),
            .in2(_gnd_net_),
            .in3(N__35397),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_15_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_15_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_13_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__35655),
            .in2(_gnd_net_),
            .in3(N__35634),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_15_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_15_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_14_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__35631),
            .in2(_gnd_net_),
            .in3(N__35613),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_15_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_15_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_15_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__35610),
            .in2(_gnd_net_),
            .in3(N__35586),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_15_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_15_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_16_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__38114),
            .in2(_gnd_net_),
            .in3(N__35583),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_15_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_15_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_17_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__35580),
            .in2(_gnd_net_),
            .in3(N__35559),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_17 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_15_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_15_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_18_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__35556),
            .in2(_gnd_net_),
            .in3(N__35538),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_15_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_19_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__35535),
            .in2(_gnd_net_),
            .in3(N__35523),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_RNO_0_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_6_LC_15_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_6_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_6_LC_15_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC841_6_LC_15_10_3  (
            .in0(N__38508),
            .in1(N__38614),
            .in2(N__38468),
            .in3(N__38259),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_15_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_15_10_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CKPA_31_LC_15_10_6  (
            .in0(N__35742),
            .in1(N__38337),
            .in2(N__43674),
            .in3(N__35673),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_11_0 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRTPU9_31_LC_15_11_0  (
            .in0(N__37976),
            .in1(N__35697),
            .in2(N__43675),
            .in3(N__43705),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31 ),
            .ltout(\delay_measurement_inst.elapsed_time_ns_1_RNIRTPU9_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_11_1 .LUT_INIT=16'b1111111100001101;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_6_LC_15_11_1  (
            .in0(N__35672),
            .in1(N__38442),
            .in2(N__35736),
            .in3(N__38262),
            .lcout(measured_delay_tr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46007),
            .ce(N__43511),
            .sr(N__45460));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_15_LC_15_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_15_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_15_LC_15_11_6 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_15_LC_15_11_6  (
            .in0(N__37953),
            .in1(N__35671),
            .in2(N__38458),
            .in3(N__35706),
            .lcout(\delay_measurement_inst.un3_elapsed_time_tr_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_15_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_15_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_15_12_0  (
            .in0(N__38546),
            .in1(N__38564),
            .in2(N__38531),
            .in3(N__38582),
            .lcout(\delay_measurement_inst.N_381 ),
            .ltout(\delay_measurement_inst.N_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_15_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_15_12_1 .LUT_INIT=16'b0001000101010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI18JP2_9_LC_15_12_1  (
            .in0(N__38451),
            .in1(N__38501),
            .in2(N__35700),
            .in3(N__38615),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_15_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_15_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIE5AP1_23_LC_15_12_2  (
            .in0(N__38817),
            .in1(N__38826),
            .in2(N__38808),
            .in3(N__38679),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_15_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_15_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_20_LC_15_12_3  (
            .in0(N__38694),
            .in1(N__35751),
            .in2(N__35691),
            .in3(N__40335),
            .lcout(\delay_measurement_inst.N_498 ),
            .ltout(\delay_measurement_inst.N_498_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_15_12_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2RFU6_7_LC_15_12_4  (
            .in0(N__38642),
            .in1(N__38663),
            .in2(N__35688),
            .in3(N__35684),
            .lcout(\delay_measurement_inst.N_384 ),
            .ltout(\delay_measurement_inst.N_384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3UDFH_6_LC_15_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3UDFH_6_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3UDFH_6_LC_15_12_5 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3UDFH_6_LC_15_12_5  (
            .in0(N__38452),
            .in1(N__35852),
            .in2(N__36000),
            .in3(N__38261),
            .lcout(\delay_measurement_inst.delay_tr_reg_5_tz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_reg_4_LC_15_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_4_LC_15_13_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_4_LC_15_13_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_4_LC_15_13_0  (
            .in0(N__38298),
            .in1(N__36388),
            .in2(N__35982),
            .in3(N__36431),
            .lcout(measured_delay_tr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \delay_measurement_inst.delay_tr_reg_5_LC_15_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_5_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_5_LC_15_13_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_5_LC_15_13_1  (
            .in0(N__36432),
            .in1(N__35926),
            .in2(N__36397),
            .in3(N__38280),
            .lcout(measured_delay_tr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_13_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_7_LC_15_13_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_7_LC_15_13_2  (
            .in0(N__38670),
            .in1(N__35858),
            .in2(N__35898),
            .in3(N__36433),
            .lcout(measured_delay_tr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_8_LC_15_13_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_8_LC_15_13_3  (
            .in0(N__36434),
            .in1(N__35823),
            .in2(N__35862),
            .in3(N__38649),
            .lcout(measured_delay_tr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \delay_measurement_inst.start_timer_hc_LC_15_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_13_4 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_15_13_4  (
            .in0(N__40719),
            .in1(N__40865),
            .in2(_gnd_net_),
            .in3(N__40759),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \delay_measurement_inst.delay_tr_reg_3_LC_15_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_3_LC_15_13_6 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_3_LC_15_13_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_3_LC_15_13_6  (
            .in0(N__38316),
            .in1(N__36387),
            .in2(N__35787),
            .in3(N__36430),
            .lcout(measured_delay_tr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \phase_controller_inst1.state_1_LC_15_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_15_13_7 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst1.state_1_LC_15_13_7  (
            .in0(N__38402),
            .in1(N__36069),
            .in2(N__36048),
            .in3(N__37932),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45989),
            .ce(),
            .sr(N__45476));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_15_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_15_14_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILDBP1_27_LC_15_14_4  (
            .in0(N__38778),
            .in1(N__38787),
            .in2(N__38769),
            .in3(N__38796),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_7_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__36064),
            .in2(_gnd_net_),
            .in3(N__36036),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_15_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_15_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_15_15_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_15_15_1  (
            .in0(N__43227),
            .in1(N__36165),
            .in2(N__36153),
            .in3(N__38230),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45974),
            .ce(),
            .sr(N__45488));
    defparam \phase_controller_inst1.state_2_LC_15_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_15_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_15_15_3 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_2_LC_15_15_3  (
            .in0(N__36150),
            .in1(N__36065),
            .in2(N__36044),
            .in3(N__36117),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45974),
            .ce(),
            .sr(N__45488));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_5 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_15_15_5  (
            .in0(N__36040),
            .in1(N__39099),
            .in2(N__40881),
            .in3(N__43165),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45974),
            .ce(),
            .sr(N__45488));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_15_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_15_7  (
            .in0(N__43396),
            .in1(N__43069),
            .in2(N__43283),
            .in3(N__36684),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45974),
            .ce(),
            .sr(N__45488));
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_15_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_15_16_0 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_7_LC_15_16_0 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_7_LC_15_16_0  (
            .in0(N__39408),
            .in1(N__46491),
            .in2(N__41238),
            .in3(N__46281),
            .lcout(measured_delay_hc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_4_LC_15_16_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_4_LC_15_16_1  (
            .in0(N__46279),
            .in1(N__41118),
            .in2(N__46499),
            .in3(N__39429),
            .lcout(measured_delay_hc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_15_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_15_16_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_30_LC_15_16_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_30_LC_15_16_2  (
            .in0(N__41321),
            .in1(N__46484),
            .in2(_gnd_net_),
            .in3(N__46278),
            .lcout(measured_delay_hc_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_15_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_5_LC_15_16_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_5_LC_15_16_3  (
            .in0(N__46280),
            .in1(N__41186),
            .in2(N__46500),
            .in3(N__42372),
            .lcout(measured_delay_hc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \phase_controller_inst1.S2_LC_15_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_15_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37945),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \delay_measurement_inst.delay_tr_reg_1_LC_15_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_1_LC_15_16_5 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_tr_reg_1_LC_15_16_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_1_LC_15_16_5  (
            .in0(N__43854),
            .in1(N__36398),
            .in2(N__36475),
            .in3(N__36440),
            .lcout(measured_delay_tr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \delay_measurement_inst.delay_tr_reg_2_LC_15_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_2_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_2_LC_15_16_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_2_LC_15_16_6  (
            .in0(N__36441),
            .in1(N__36349),
            .in2(N__36402),
            .in3(N__38367),
            .lcout(measured_delay_tr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_16_7 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_15_16_7  (
            .in0(N__37838),
            .in1(N__40837),
            .in2(_gnd_net_),
            .in3(N__39847),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45970),
            .ce(),
            .sr(N__45492));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__36663),
            .in2(N__36333),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_2_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__36312),
            .in2(_gnd_net_),
            .in3(N__36282),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_3_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__36279),
            .in2(N__36261),
            .in3(N__36234),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_4_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__36231),
            .in2(_gnd_net_),
            .in3(N__36201),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_5_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__36198),
            .in2(_gnd_net_),
            .in3(N__36168),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_6_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__36636),
            .in2(_gnd_net_),
            .in3(N__36606),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_7_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__38870),
            .in2(_gnd_net_),
            .in3(N__36603),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_8_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__38843),
            .in2(_gnd_net_),
            .in3(N__36600),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_9_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__36864),
            .in2(_gnd_net_),
            .in3(N__36597),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_10_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__36593),
            .in2(_gnd_net_),
            .in3(N__36573),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_11_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__36569),
            .in2(_gnd_net_),
            .in3(N__36549),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_12_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__36545),
            .in2(_gnd_net_),
            .in3(N__36525),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_13_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__36522),
            .in2(_gnd_net_),
            .in3(N__36492),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_14_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__36749),
            .in2(_gnd_net_),
            .in3(N__36729),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_15_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__36725),
            .in2(_gnd_net_),
            .in3(N__36705),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_16_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__36701),
            .in2(_gnd_net_),
            .in3(N__36675),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_17_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__36885),
            .in2(_gnd_net_),
            .in3(N__36672),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_18_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__36843),
            .in2(_gnd_net_),
            .in3(N__36669),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_RNO_0_19_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__36648),
            .in2(_gnd_net_),
            .in3(N__36666),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__39078),
            .in2(_gnd_net_),
            .in3(N__43155),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_20_0 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_20_0  (
            .in0(N__43110),
            .in1(N__43453),
            .in2(N__43336),
            .in3(N__36654),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45951),
            .ce(),
            .sr(N__45524));
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_15_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_10_LC_15_20_1 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_10_LC_15_20_1  (
            .in0(N__46439),
            .in1(N__39219),
            .in2(N__41075),
            .in3(N__46255),
            .lcout(measured_delay_hc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45951),
            .ce(),
            .sr(N__45524));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_20_2 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_20_2  (
            .in0(N__43108),
            .in1(N__43452),
            .in2(N__43334),
            .in3(N__36891),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45951),
            .ce(),
            .sr(N__45524));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_20_3 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_20_3  (
            .in0(N__43451),
            .in1(N__36873),
            .in2(N__43126),
            .in3(N__43311),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45951),
            .ce(),
            .sr(N__45524));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_20_6 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_20_6  (
            .in0(N__43109),
            .in1(N__36849),
            .in2(N__43335),
            .in3(N__43454),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45951),
            .ce(),
            .sr(N__45524));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_15_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_15_21_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__46730),
            .in2(_gnd_net_),
            .in3(N__47021),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45949),
            .ce(N__38937),
            .sr(N__45533));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_15_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_15_21_2 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_15_21_2  (
            .in0(N__46731),
            .in1(N__46995),
            .in2(_gnd_net_),
            .in3(N__46830),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45949),
            .ce(N__38937),
            .sr(N__45533));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_15_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_15_21_5 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_15_21_5  (
            .in0(N__46828),
            .in1(N__46732),
            .in2(_gnd_net_),
            .in3(N__46643),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45949),
            .ce(N__38937),
            .sr(N__45533));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_15_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_15_21_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_15_21_7  (
            .in0(N__46829),
            .in1(N__46733),
            .in2(_gnd_net_),
            .in3(N__41868),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45949),
            .ce(N__38937),
            .sr(N__45533));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_22_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__36795),
            .in2(N__37118),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__36774),
            .in2(N__37091),
            .in3(N__36753),
            .lcout(\delay_measurement_inst.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__37061),
            .in2(N__37119),
            .in3(N__37095),
            .lcout(\delay_measurement_inst.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__37037),
            .in2(N__37092),
            .in3(N__37065),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__37062),
            .in2(N__37013),
            .in3(N__37041),
            .lcout(\delay_measurement_inst.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__37038),
            .in2(N__36983),
            .in3(N__37017),
            .lcout(\delay_measurement_inst.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__36953),
            .in2(N__37014),
            .in3(N__36987),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(N__36921),
            .in2(N__36984),
            .in3(N__36957),
            .lcout(\delay_measurement_inst.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__45946),
            .ce(N__37860),
            .sr(N__45540));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(N__36954),
            .in2(N__37364),
            .in3(N__36924),
            .lcout(\delay_measurement_inst.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(N__36920),
            .in2(N__37337),
            .in3(N__36894),
            .lcout(\delay_measurement_inst.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_23_2  (
            .in0(_gnd_net_),
            .in1(N__37307),
            .in2(N__37365),
            .in3(N__37341),
            .lcout(\delay_measurement_inst.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__37286),
            .in2(N__37338),
            .in3(N__37311),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_23_4  (
            .in0(_gnd_net_),
            .in1(N__37308),
            .in2(N__37262),
            .in3(N__37290),
            .lcout(\delay_measurement_inst.delay_hc_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_23_5  (
            .in0(_gnd_net_),
            .in1(N__37287),
            .in2(N__37232),
            .in3(N__37266),
            .lcout(\delay_measurement_inst.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_23_6  (
            .in0(_gnd_net_),
            .in1(N__37203),
            .in2(N__37263),
            .in3(N__37236),
            .lcout(\delay_measurement_inst.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_23_7  (
            .in0(_gnd_net_),
            .in1(N__37173),
            .in2(N__37233),
            .in3(N__37206),
            .lcout(\delay_measurement_inst.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__45943),
            .ce(N__37859),
            .sr(N__45546));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_24_0  (
            .in0(_gnd_net_),
            .in1(N__37202),
            .in2(N__37142),
            .in3(N__37176),
            .lcout(\delay_measurement_inst.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__37172),
            .in2(N__37607),
            .in3(N__37146),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__37577),
            .in2(N__37143),
            .in3(N__37611),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_24_3  (
            .in0(_gnd_net_),
            .in1(N__37553),
            .in2(N__37608),
            .in3(N__37581),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__37578),
            .in2(N__37529),
            .in3(N__37557),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_24_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__37554),
            .in2(N__37499),
            .in3(N__37533),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_24_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_24_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_24_6  (
            .in0(_gnd_net_),
            .in1(N__37470),
            .in2(N__37530),
            .in3(N__37503),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_24_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_24_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_24_7  (
            .in0(_gnd_net_),
            .in1(N__37440),
            .in2(N__37500),
            .in3(N__37473),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__45939),
            .ce(N__37858),
            .sr(N__45554));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_25_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__37469),
            .in2(N__37391),
            .in3(N__37443),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__45935),
            .ce(N__37857),
            .sr(N__45559));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_25_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_25_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_25_1  (
            .in0(_gnd_net_),
            .in1(N__37439),
            .in2(N__37889),
            .in3(N__37413),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__45935),
            .ce(N__37857),
            .sr(N__45559));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_25_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_25_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__37410),
            .in2(N__37392),
            .in3(N__37368),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__45935),
            .ce(N__37857),
            .sr(N__45559));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_25_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_25_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_25_3  (
            .in0(_gnd_net_),
            .in1(N__37908),
            .in2(N__37890),
            .in3(N__37866),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__45935),
            .ce(N__37857),
            .sr(N__45559));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_25_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_25_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_25_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37863),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45935),
            .ce(N__37857),
            .sr(N__45559));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_26_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_26_1 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_26_1  (
            .in0(N__37839),
            .in1(N__40842),
            .in2(_gnd_net_),
            .in3(N__39864),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_462_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_27_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_27_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_27_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_27_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39863),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_5_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_5_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39788),
            .lcout(\delay_measurement_inst.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46060),
            .ce(N__43825),
            .sr(N__45440));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI104I_2_LC_16_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI104I_2_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI104I_2_LC_16_6_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI104I_2_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__38509),
            .in2(_gnd_net_),
            .in3(N__38356),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_16_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_16_7_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_16_7_1  (
            .in0(N__42849),
            .in1(N__42629),
            .in2(_gnd_net_),
            .in3(N__42793),
            .lcout(\phase_controller_inst1.stoper_tr.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37653),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNI7NN7_0_LC_16_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.state_RNI7NN7_0_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__38095),
            .in2(_gnd_net_),
            .in3(N__38084),
            .lcout(\phase_controller_inst1.state_RNI7NN7Z0Z_0 ),
            .ltout(\phase_controller_inst1.state_RNI7NN7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_16_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_16_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_16_8_1 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_16_8_1  (
            .in0(N__38376),
            .in1(N__42918),
            .in2(N__38235),
            .in3(N__38232),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46044),
            .ce(),
            .sr(N__45443));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_16_8_3 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_16_8_3  (
            .in0(N__38099),
            .in1(N__38160),
            .in2(N__38133),
            .in3(N__42681),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46044),
            .ce(),
            .sr(N__45443));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_8_4 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_16_8_4  (
            .in0(N__42628),
            .in1(N__42812),
            .in2(N__42954),
            .in3(N__38124),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46044),
            .ce(),
            .sr(N__45443));
    defparam \phase_controller_inst1.state_0_LC_16_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_16_8_5 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst1.state_0_LC_16_8_5  (
            .in0(N__38085),
            .in1(N__37947),
            .in2(N__38100),
            .in3(N__38401),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46044),
            .ce(),
            .sr(N__45443));
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_16_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_16_LC_16_9_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_16_LC_16_9_1  (
            .in0(N__43721),
            .in1(N__43647),
            .in2(_gnd_net_),
            .in3(N__38751),
            .lcout(measured_delay_tr_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46036),
            .ce(N__43521),
            .sr(N__45446));
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_9_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_9_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_19_LC_16_9_7  (
            .in0(N__43722),
            .in1(N__43648),
            .in2(_gnd_net_),
            .in3(N__38720),
            .lcout(measured_delay_tr_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46036),
            .ce(N__43521),
            .sr(N__45446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_10_0  (
            .in0(N__38750),
            .in1(N__38719),
            .in2(N__43806),
            .in3(N__43577),
            .lcout(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16 ),
            .ltout(\delay_measurement_inst.elapsed_time_ns_1_RNIM96P1_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH1A23_1_LC_16_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH1A23_1_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH1A23_1_LC_16_10_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH1A23_1_LC_16_10_1  (
            .in0(N__38331),
            .in1(N__38322),
            .in2(N__37965),
            .in3(N__37962),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__37946),
            .in2(_gnd_net_),
            .in3(N__38403),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICA841_2_LC_16_10_3  (
            .in0(N__43576),
            .in1(N__38311),
            .in2(N__38721),
            .in3(N__38363),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_10_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIOKG82_16_LC_16_10_4  (
            .in0(N__43801),
            .in1(N__38749),
            .in2(N__38340),
            .in3(N__38330),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__38276),
            .in2(_gnd_net_),
            .in3(N__38294),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_373_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_16_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_16_10_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7GAF_1_LC_16_10_7  (
            .in0(N__38613),
            .in1(N__38312),
            .in2(N__43850),
            .in3(N__38260),
            .lcout(\delay_measurement_inst.delay_tr_timer.un3_elapsed_time_tr_0_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__43881),
            .in2(N__39758),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__39731),
            .in2(N__39795),
            .in3(N__38283),
            .lcout(\delay_measurement_inst.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__39710),
            .in2(N__39759),
            .in3(N__38265),
            .lcout(\delay_measurement_inst.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__39732),
            .in2(N__39681),
            .in3(N__38238),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__40079),
            .in2(N__39711),
            .in3(N__38652),
            .lcout(\delay_measurement_inst.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__39677),
            .in2(N__40058),
            .in3(N__38631),
            .lcout(\delay_measurement_inst.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__40080),
            .in2(N__40028),
            .in3(N__38592),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__39991),
            .in2(N__40059),
            .in3(N__38571),
            .lcout(\delay_measurement_inst.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__46017),
            .ce(N__43826),
            .sr(N__45457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__40029),
            .in2(N__39965),
            .in3(N__38553),
            .lcout(\delay_measurement_inst.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__39938),
            .in2(N__39999),
            .in3(N__38535),
            .lcout(\delay_measurement_inst.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__39917),
            .in2(N__39966),
            .in3(N__38514),
            .lcout(\delay_measurement_inst.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__39939),
            .in2(N__39894),
            .in3(N__38472),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__39918),
            .in2(N__40325),
            .in3(N__38754),
            .lcout(\delay_measurement_inst.delay_tr_reg3lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__39890),
            .in2(N__40295),
            .in3(N__38730),
            .lcout(\delay_measurement_inst.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__40268),
            .in2(N__40326),
            .in3(N__38727),
            .lcout(\delay_measurement_inst.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__40232),
            .in2(N__40296),
            .in3(N__38724),
            .lcout(\delay_measurement_inst.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__46008),
            .ce(N__43827),
            .sr(N__45461));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__40269),
            .in2(N__40208),
            .in3(N__38697),
            .lcout(\delay_measurement_inst.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__40236),
            .in2(N__40181),
            .in3(N__38688),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__40151),
            .in2(N__40209),
            .in3(N__38685),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__40121),
            .in2(N__40182),
            .in3(N__38682),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__40100),
            .in2(N__40152),
            .in3(N__38673),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__40122),
            .in2(N__40691),
            .in3(N__38820),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__40101),
            .in2(N__40664),
            .in3(N__38811),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__40628),
            .in2(N__40692),
            .in3(N__38799),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__45999),
            .ce(N__43829),
            .sr(N__45468));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__40665),
            .in2(N__40601),
            .in3(N__38790),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__45990),
            .ce(N__43830),
            .sr(N__45477));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__40574),
            .in2(N__40635),
            .in3(N__38781),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__45990),
            .ce(N__43830),
            .sr(N__45477));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__40554),
            .in2(N__40602),
            .in3(N__38772),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__45990),
            .ce(N__43830),
            .sr(N__45477));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__40575),
            .in2(N__40407),
            .in3(N__38760),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_trZ0Z_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__45990),
            .ce(N__43830),
            .sr(N__45477));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38757),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45990),
            .ce(N__43830),
            .sr(N__45477));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_15_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_0_LC_16_15_0  (
            .in0(N__43046),
            .in1(N__43428),
            .in2(N__43284),
            .in3(N__43172),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45980),
            .ce(N__42502),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.hc_state_0_LC_16_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.hc_state_0_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.hc_state_0_LC_16_15_2 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \delay_measurement_inst.hc_state_0_LC_16_15_2  (
            .in0(N__40708),
            .in1(N__40858),
            .in2(_gnd_net_),
            .in3(N__40760),
            .lcout(\delay_measurement_inst.hc_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45980),
            .ce(N__42502),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_3_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_3_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_3_LC_16_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_3_LC_16_17_5  (
            .in0(N__41644),
            .in1(N__46131),
            .in2(N__41187),
            .in3(N__41934),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_LC_16_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_LC_16_17_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_1_0_a3_0_LC_16_17_6  (
            .in0(N__41224),
            .in1(N__41097),
            .in2(N__38889),
            .in3(N__42076),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.N_316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_i_LC_16_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_i_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto8_i_LC_16_17_7 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto8_i_LC_16_17_7  (
            .in0(N__40946),
            .in1(N__41293),
            .in2(N__38886),
            .in3(N__41225),
            .lcout(\phase_controller_inst1.stoper_hc.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_16_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_16_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_16_18_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_16_18_0  (
            .in0(N__43071),
            .in1(N__43315),
            .in2(N__38883),
            .in3(N__43443),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45965),
            .ce(),
            .sr(N__45499));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_16_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_16_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_16_18_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_16_18_1  (
            .in0(N__43442),
            .in1(N__43072),
            .in2(N__43337),
            .in3(N__38853),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45965),
            .ce(),
            .sr(N__45499));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_2_0_a2_LC_16_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_2_0_a2_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto13_2_0_a2_LC_16_18_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto13_2_0_a2_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__40970),
            .in2(_gnd_net_),
            .in3(N__41018),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un2_startlt31_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3_2_LC_16_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3_2_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3_2_LC_16_18_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3_2_LC_16_18_4  (
            .in0(N__41070),
            .in1(N__41828),
            .in2(N__38829),
            .in3(N__42259),
            .lcout(\phase_controller_inst1.stoper_hc.un1_startlto19_3_i_a3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_16_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_11_LC_16_18_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_11_LC_16_18_6  (
            .in0(N__39258),
            .in1(N__46461),
            .in2(N__41029),
            .in3(N__46265),
            .lcout(measured_delay_hc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45965),
            .ce(),
            .sr(N__45499));
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_16_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_16_18_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_12_LC_16_18_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_12_LC_16_18_7  (
            .in0(N__46266),
            .in1(N__40971),
            .in2(N__46494),
            .in3(N__39276),
            .lcout(measured_delay_hc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45965),
            .ce(),
            .sr(N__45499));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_16_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_16_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_16_19_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_16_19_0  (
            .in0(N__41456),
            .in1(N__46130),
            .in2(N__41769),
            .in3(N__46914),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_16_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_16_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_16_19_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_16_19_1  (
            .in0(N__46912),
            .in1(N__41746),
            .in2(N__41500),
            .in3(N__41241),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_16_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_16_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_16_19_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_16_19_2  (
            .in0(N__41455),
            .in1(N__42261),
            .in2(N__41768),
            .in3(N__46913),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_19_3 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_16_19_3  (
            .in0(N__46909),
            .in1(N__46746),
            .in2(N__41595),
            .in3(N__41458),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_16_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_16_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_16_19_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_16_19_4  (
            .in0(N__41457),
            .in1(N__41191),
            .in2(N__41770),
            .in3(N__46915),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_16_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_16_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_16_19_5 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_16_19_5  (
            .in0(N__46911),
            .in1(N__46747),
            .in2(N__41295),
            .in3(N__41460),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_16_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_16_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_16_19_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_16_19_7  (
            .in0(N__46910),
            .in1(N__41646),
            .in2(N__41655),
            .in3(N__41459),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45959),
            .ce(N__38933),
            .sr(N__45508));
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_0_LC_16_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_0_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_0_LC_16_20_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_i_0_LC_16_20_0  (
            .in0(N__41669),
            .in1(N__39108),
            .in2(N__42005),
            .in3(N__46702),
            .lcout(\phase_controller_inst1.stoper_hc.un3_start_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_o2_1_LC_16_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_o2_1_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_o2_1_LC_16_20_2 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_o2_1_LC_16_20_2  (
            .in0(N__41935),
            .in1(N__41637),
            .in2(_gnd_net_),
            .in3(N__46129),
            .lcout(\phase_controller_inst1.stoper_hc.N_406 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_1_LC_16_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_1_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_1_LC_16_20_3 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_1_LC_16_20_3  (
            .in0(N__46701),
            .in1(N__41668),
            .in2(N__39102),
            .in3(N__47020),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_16_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_16_20_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_RNILRMG_0_LC_16_20_4  (
            .in0(_gnd_net_),
            .in1(N__43070),
            .in2(_gnd_net_),
            .in3(N__43397),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_8_LC_16_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_8_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_8_LC_16_20_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_8_LC_16_20_5  (
            .in0(N__41282),
            .in1(N__41028),
            .in2(N__40990),
            .in3(N__41239),
            .lcout(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_7_LC_16_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_7_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_7_LC_16_20_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_7_LC_16_20_6  (
            .in0(N__41867),
            .in1(N__41373),
            .in2(N__41593),
            .in3(N__41119),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_LC_16_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_LC_16_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_LC_16_20_7  (
            .in0(N__39060),
            .in1(N__39051),
            .in2(N__39054),
            .in3(N__39045),
            .lcout(\phase_controller_inst1.stoper_hc.N_459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_5_LC_16_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_5_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_5_LC_16_21_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_5_LC_16_21_0  (
            .in0(N__42257),
            .in1(N__46637),
            .in2(_gnd_net_),
            .in3(N__46983),
            .lcout(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3_18_LC_16_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3_18_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3_18_LC_16_21_1 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3_18_LC_16_21_1  (
            .in0(N__41582),
            .in1(N__39282),
            .in2(_gnd_net_),
            .in3(N__42258),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_3Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_6_LC_16_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_6_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_6_LC_16_21_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_start_i_a2_0_6_LC_16_21_4  (
            .in0(N__41069),
            .in1(N__40938),
            .in2(N__41827),
            .in3(N__41195),
            .lcout(\phase_controller_inst1.stoper_hc.un3_start_i_a2_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_19_LC_16_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_19_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_19_LC_16_21_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_19_LC_16_21_7  (
            .in0(_gnd_net_),
            .in1(N__41990),
            .in2(_gnd_net_),
            .in3(N__46791),
            .lcout(\phase_controller_inst1.stoper_hc.N_453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2_18_LC_16_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2_18_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2_18_LC_16_22_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2_18_LC_16_22_0  (
            .in0(N__41859),
            .in1(N__46642),
            .in2(N__41998),
            .in3(N__46982),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_2Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_16_LC_16_22_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_16_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_16_LC_16_22_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TRB1_16_LC_16_22_2  (
            .in0(N__41953),
            .in1(N__39424),
            .in2(N__39464),
            .in3(N__42358),
            .lcout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_22_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIDD01_10_LC_16_22_3  (
            .in0(N__39269),
            .in1(N__39251),
            .in2(N__39236),
            .in3(N__39215),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7_19_LC_16_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7_19_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7_19_LC_16_22_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7_19_LC_16_22_4  (
            .in0(N__39204),
            .in1(N__46515),
            .in2(N__39486),
            .in3(N__39189),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_7Z0Z_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_19_LC_16_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_19_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_19_LC_16_22_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_19_LC_16_22_5  (
            .in0(N__41304),
            .in1(N__39174),
            .in2(N__39159),
            .in3(N__39540),
            .lcout(\phase_controller_inst1.stoper_hc.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_22_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIA6E01_16_LC_16_22_6  (
            .in0(N__41954),
            .in1(N__41884),
            .in2(N__42044),
            .in3(N__39460),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_o2_0_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_14_LC_16_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_14_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_14_LC_16_23_1 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_14_LC_16_23_1  (
            .in0(N__39155),
            .in1(N__39137),
            .in2(_gnd_net_),
            .in3(N__39307),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGMFO5_15_LC_16_23_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGMFO5_15_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGMFO5_15_LC_16_23_2 .LUT_INIT=16'b1100110001000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGMFO5_15_LC_16_23_2  (
            .in0(N__42278),
            .in1(N__39294),
            .in2(N__39120),
            .in3(N__39117),
            .lcout(\delay_measurement_inst.N_332 ),
            .ltout(\delay_measurement_inst.N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICFUBH_31_LC_16_23_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICFUBH_31_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICFUBH_31_LC_16_23_3 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICFUBH_31_LC_16_23_3  (
            .in0(N__39651),
            .in1(N__39363),
            .in2(N__39111),
            .in3(N__42306),
            .lcout(\delay_measurement_inst.N_298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_23_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_23_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_4_LC_16_23_4  (
            .in0(N__42277),
            .in1(N__39523),
            .in2(N__39404),
            .in3(N__39425),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHVTL_7_LC_16_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHVTL_7_LC_16_23_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHVTL_7_LC_16_23_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHVTL_7_LC_16_23_5  (
            .in0(_gnd_net_),
            .in1(N__39397),
            .in2(_gnd_net_),
            .in3(N__42276),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_318_1 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_318_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO11I2_18_LC_16_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO11I2_18_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO11I2_18_LC_16_23_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIO11I2_18_LC_16_23_6  (
            .in0(N__42040),
            .in1(N__41885),
            .in2(N__39384),
            .in3(N__39381),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un1_elapsed_time_hc_1_i_a3_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_14_LC_16_23_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_14_LC_16_23_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_14_LC_16_23_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8MV5_14_LC_16_23_7  (
            .in0(N__39375),
            .in1(N__39503),
            .in2(N__39366),
            .in3(N__39308),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_16_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_16_24_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_16_24_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRQ8G_21_LC_16_24_0  (
            .in0(N__39357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39351),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_24_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_24_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_24_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2JIP2_20_LC_16_24_1  (
            .in0(N__39345),
            .in1(N__39564),
            .in2(N__39336),
            .in3(N__39597),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_328 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOFS27_1_LC_16_24_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOFS27_1_LC_16_24_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOFS27_1_LC_16_24_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOFS27_1_LC_16_24_2  (
            .in0(N__39315),
            .in1(N__42345),
            .in2(N__39333),
            .in3(N__39330),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI71JB5_6_LC_16_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI71JB5_6_LC_16_24_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI71JB5_6_LC_16_24_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI71JB5_6_LC_16_24_5  (
            .in0(N__39321),
            .in1(N__39314),
            .in2(N__39504),
            .in3(N__39293),
            .lcout(\delay_measurement_inst.N_318 ),
            .ltout(\delay_measurement_inst.N_318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDM4FI_31_LC_16_24_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDM4FI_31_LC_16_24_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDM4FI_31_LC_16_24_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDM4FI_31_LC_16_24_6  (
            .in0(N__39647),
            .in1(N__39633),
            .in2(N__39627),
            .in3(N__42318),
            .lcout(\delay_measurement_inst.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_16_24_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_16_24_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_16_24_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_16_24_7  (
            .in0(N__39624),
            .in1(N__39618),
            .in2(N__39612),
            .in3(N__39603),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_25_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_25_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_25_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_16_25_0  (
            .in0(N__39591),
            .in1(N__39585),
            .in2(N__39579),
            .in3(N__39570),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg_3_i_a2_1_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0_19_LC_16_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0_19_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0_19_LC_16_25_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0_19_LC_16_25_3  (
            .in0(_gnd_net_),
            .in1(N__39558),
            .in2(_gnd_net_),
            .in3(N__39440),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_0Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI21LR_6_LC_16_25_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI21LR_6_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI21LR_6_LC_16_25_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI21LR_6_LC_16_25_4  (
            .in0(_gnd_net_),
            .in1(N__39531),
            .in2(_gnd_net_),
            .in3(N__42335),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_408 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_16_26_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_16_26_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_26_LC_16_26_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_26_LC_16_26_1  (
            .in0(N__39479),
            .in1(N__46380),
            .in2(_gnd_net_),
            .in3(N__46222),
            .lcout(measured_delay_hc_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45936),
            .ce(),
            .sr(N__45560));
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_16_26_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_16_26_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_17_LC_16_26_3 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_17_LC_16_26_3  (
            .in0(N__39465),
            .in1(N__46378),
            .in2(N__46641),
            .in3(N__46220),
            .lcout(measured_delay_hc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45936),
            .ce(),
            .sr(N__45560));
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_16_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_16_26_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_20_LC_16_26_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_20_LC_16_26_5  (
            .in0(N__39441),
            .in1(N__46379),
            .in2(_gnd_net_),
            .in3(N__46221),
            .lcout(measured_delay_hc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45936),
            .ce(),
            .sr(N__45560));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_28_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_28_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_16_28_2  (
            .in0(_gnd_net_),
            .in1(N__40838),
            .in2(_gnd_net_),
            .in3(N__39856),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_461_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC1_LC_17_6_7.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC1_LC_17_6_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC1_LC_17_6_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC1_LC_17_6_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39813),
            .lcout(delay_hc_d1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46061),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_DELAY_HC2_LC_17_7_4.C_ON=1'b0;
    defparam SB_DFF_inst_DELAY_HC2_LC_17_7_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_DELAY_HC2_LC_17_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_DELAY_HC2_LC_17_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39804),
            .lcout(delay_hc_d2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46058),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_8_0  (
            .in0(N__40461),
            .in1(N__43870),
            .in2(_gnd_net_),
            .in3(N__39798),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_8_1  (
            .in0(N__40456),
            .in1(N__39781),
            .in2(_gnd_net_),
            .in3(N__39762),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_8_2  (
            .in0(N__40462),
            .in1(N__39751),
            .in2(_gnd_net_),
            .in3(N__39735),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_8_3  (
            .in0(N__40457),
            .in1(N__39730),
            .in2(_gnd_net_),
            .in3(N__39714),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_8_4  (
            .in0(N__40463),
            .in1(N__39703),
            .in2(_gnd_net_),
            .in3(N__39684),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_8_5  (
            .in0(N__40458),
            .in1(N__39673),
            .in2(_gnd_net_),
            .in3(N__39654),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_8_6  (
            .in0(N__40460),
            .in1(N__40078),
            .in2(_gnd_net_),
            .in3(N__40062),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_8_7  (
            .in0(N__40459),
            .in1(N__40046),
            .in2(_gnd_net_),
            .in3(N__40032),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__46053),
            .ce(N__40385),
            .sr(N__45441));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_9_0  (
            .in0(N__40525),
            .in1(N__40021),
            .in2(_gnd_net_),
            .in3(N__40002),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_9_1  (
            .in0(N__40529),
            .in1(N__39995),
            .in2(_gnd_net_),
            .in3(N__39969),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_9_2  (
            .in0(N__40522),
            .in1(N__39958),
            .in2(_gnd_net_),
            .in3(N__39942),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_9_3  (
            .in0(N__40526),
            .in1(N__39937),
            .in2(_gnd_net_),
            .in3(N__39921),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_9_4  (
            .in0(N__40523),
            .in1(N__39911),
            .in2(_gnd_net_),
            .in3(N__39897),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_9_5  (
            .in0(N__40527),
            .in1(N__39886),
            .in2(_gnd_net_),
            .in3(N__39867),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_9_6  (
            .in0(N__40524),
            .in1(N__40313),
            .in2(_gnd_net_),
            .in3(N__40299),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_9_7  (
            .in0(N__40528),
            .in1(N__40288),
            .in2(_gnd_net_),
            .in3(N__40272),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__46045),
            .ce(N__40377),
            .sr(N__45444));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_10_0  (
            .in0(N__40530),
            .in1(N__40258),
            .in2(_gnd_net_),
            .in3(N__40239),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_10_1  (
            .in0(N__40485),
            .in1(N__40231),
            .in2(_gnd_net_),
            .in3(N__40212),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_10_2  (
            .in0(N__40531),
            .in1(N__40201),
            .in2(_gnd_net_),
            .in3(N__40185),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_10_3  (
            .in0(N__40486),
            .in1(N__40169),
            .in2(_gnd_net_),
            .in3(N__40155),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_10_4  (
            .in0(N__40532),
            .in1(N__40144),
            .in2(_gnd_net_),
            .in3(N__40125),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_10_5  (
            .in0(N__40487),
            .in1(N__40120),
            .in2(_gnd_net_),
            .in3(N__40104),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_10_6  (
            .in0(N__40533),
            .in1(N__40099),
            .in2(_gnd_net_),
            .in3(N__40083),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_10_7  (
            .in0(N__40488),
            .in1(N__40684),
            .in2(_gnd_net_),
            .in3(N__40668),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__46037),
            .ce(N__40386),
            .sr(N__45447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_11_0  (
            .in0(N__40489),
            .in1(N__40657),
            .in2(_gnd_net_),
            .in3(N__40638),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__46026),
            .ce(N__40378),
            .sr(N__45455));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_11_1  (
            .in0(N__40493),
            .in1(N__40627),
            .in2(_gnd_net_),
            .in3(N__40605),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__46026),
            .ce(N__40378),
            .sr(N__45455));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_11_2  (
            .in0(N__40490),
            .in1(N__40594),
            .in2(_gnd_net_),
            .in3(N__40578),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__46026),
            .ce(N__40378),
            .sr(N__45455));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_11_3  (
            .in0(N__40494),
            .in1(N__40573),
            .in2(_gnd_net_),
            .in3(N__40557),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__46026),
            .ce(N__40378),
            .sr(N__45455));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_11_4  (
            .in0(N__40491),
            .in1(N__40550),
            .in2(_gnd_net_),
            .in3(N__40536),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__46026),
            .ce(N__40378),
            .sr(N__45455));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_11_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_11_5  (
            .in0(N__40400),
            .in1(N__40492),
            .in2(_gnd_net_),
            .in3(N__40410),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46026),
            .ce(N__40378),
            .sr(N__45455));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_17_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_17_12_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__40347),
            .in2(_gnd_net_),
            .in3(N__40341),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_reg_5_i_o2_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_17_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_17_13_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_17_13_4  (
            .in0(N__43286),
            .in1(N__42996),
            .in2(_gnd_net_),
            .in3(N__43401),
            .lcout(\phase_controller_inst1.stoper_hc.time_passed_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_17_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_17_13_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.stop_timer_hc_LC_17_13_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_17_13_7  (
            .in0(N__40715),
            .in1(N__40866),
            .in2(N__45624),
            .in3(N__40749),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46009),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_17_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_17_14_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_17_14_4  (
            .in0(N__44584),
            .in1(N__44429),
            .in2(_gnd_net_),
            .in3(N__44300),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_hc.time_passed_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_17_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_17_14_5 .LUT_INIT=16'b1010100010101100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_17_14_5  (
            .in0(N__40782),
            .in1(N__43944),
            .in2(N__40797),
            .in3(N__47070),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46000),
            .ce(),
            .sr(N__45469));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_17_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_17_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNINF2L_0_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__44428),
            .in2(_gnd_net_),
            .in3(N__44299),
            .lcout(\phase_controller_inst2.stoper_hc.time_passed11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_14_7 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_14_7  (
            .in0(N__44301),
            .in1(N__44585),
            .in2(N__44474),
            .in3(N__43998),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46000),
            .ce(),
            .sr(N__45469));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_1 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_1  (
            .in0(N__44476),
            .in1(N__44338),
            .in2(N__44641),
            .in3(N__43962),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45991),
            .ce(),
            .sr(N__45478));
    defparam \delay_measurement_inst.prev_hc_sig_LC_17_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.prev_hc_sig_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.prev_hc_sig_LC_17_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.prev_hc_sig_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40761),
            .lcout(\delay_measurement_inst.prev_hc_sigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45991),
            .ce(),
            .sr(N__45478));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_3 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_3  (
            .in0(N__44477),
            .in1(N__44019),
            .in2(N__44642),
            .in3(N__44339),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45991),
            .ce(),
            .sr(N__45478));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_7  (
            .in0(N__44475),
            .in1(N__44337),
            .in2(N__44640),
            .in3(N__43971),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45991),
            .ce(),
            .sr(N__45478));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_16_1 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_16_1  (
            .in0(N__43896),
            .in1(N__44482),
            .in2(N__44663),
            .in3(N__44345),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45981),
            .ce(),
            .sr(N__45484));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_2 .LUT_INIT=16'b1100100010001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_2  (
            .in0(N__44342),
            .in1(N__44085),
            .in2(N__44507),
            .in3(N__44639),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45981),
            .ce(),
            .sr(N__45484));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_4  (
            .in0(N__44341),
            .in1(N__44632),
            .in2(N__44506),
            .in3(N__44094),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45981),
            .ce(),
            .sr(N__45484));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_16_5 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_16_5  (
            .in0(N__43986),
            .in1(N__44481),
            .in2(N__44662),
            .in3(N__44344),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45981),
            .ce(),
            .sr(N__45484));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_7 .LUT_INIT=16'b1110110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_7  (
            .in0(N__44631),
            .in1(N__44343),
            .in2(N__44505),
            .in3(N__44073),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45981),
            .ce(),
            .sr(N__45484));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_17_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_17_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_17_17_0 .LUT_INIT=16'b0000101100001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_17_17_0  (
            .in0(N__41294),
            .in1(N__41464),
            .in2(N__46755),
            .in3(N__46939),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45975),
            .ce(N__46561),
            .sr(N__45489));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_17_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_17_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_17_17_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_17_17_1  (
            .in0(N__46937),
            .in1(N__41778),
            .in2(N__41497),
            .in3(N__40950),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45975),
            .ce(N__46561),
            .sr(N__45489));
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_17_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_17_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_0_LC_17_17_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_0_LC_17_17_4  (
            .in0(N__42077),
            .in1(N__41463),
            .in2(N__41780),
            .in3(N__46938),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45975),
            .ce(N__46561),
            .sr(N__45489));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_17_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_17_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_17_17_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_17_17_5  (
            .in0(N__46935),
            .in1(N__41936),
            .in2(N__41495),
            .in3(N__40898),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45975),
            .ce(N__46561),
            .sr(N__45489));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_17_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_17_17_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_17_17_6  (
            .in0(N__41240),
            .in1(N__41465),
            .in2(N__41781),
            .in3(N__46940),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45975),
            .ce(N__46561),
            .sr(N__45489));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_17_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_17_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_17_17_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_17_17_7  (
            .in0(N__46936),
            .in1(N__41771),
            .in2(N__41496),
            .in3(N__41196),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45975),
            .ce(N__46561),
            .sr(N__45489));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_18_LC_17_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_18_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_18_LC_17_18_1 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_o2_18_LC_17_18_1  (
            .in0(N__41375),
            .in1(N__41151),
            .in2(N__41142),
            .in3(N__41133),
            .lcout(\phase_controller_inst1.stoper_hc.N_405 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_405_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_17_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_17_18_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_17_18_2  (
            .in0(N__46890),
            .in1(N__41764),
            .in2(N__41127),
            .in3(N__46128),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45971),
            .ce(N__46579),
            .sr(N__45493));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_17_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_17_18_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_17_18_3  (
            .in0(N__41124),
            .in1(N__41462),
            .in2(N__41779),
            .in3(N__46892),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45971),
            .ce(N__46579),
            .sr(N__45493));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_17_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_17_18_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_17_18_7  (
            .in0(N__41763),
            .in1(N__41461),
            .in2(N__41079),
            .in3(N__46891),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45971),
            .ce(N__46579),
            .sr(N__45493));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_17_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_17_19_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_17_19_0  (
            .in0(N__41733),
            .in1(N__41475),
            .in2(N__41030),
            .in3(N__46835),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45966),
            .ce(N__46577),
            .sr(N__45500));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_17_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_17_19_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_17_19_1  (
            .in0(N__46833),
            .in1(N__42260),
            .in2(N__41499),
            .in3(N__41736),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45966),
            .ce(N__46577),
            .sr(N__45500));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_17_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_17_19_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_17_19_2  (
            .in0(N__41734),
            .in1(N__41476),
            .in2(N__40992),
            .in3(N__46836),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45966),
            .ce(N__46577),
            .sr(N__45500));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_17_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_17_19_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_17_19_3  (
            .in0(N__46832),
            .in1(N__41829),
            .in2(N__41498),
            .in3(N__41735),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45966),
            .ce(N__46577),
            .sr(N__45500));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_3_LC_17_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_3_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_3_LC_17_19_6 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_0_0_3_LC_17_19_6  (
            .in0(N__41670),
            .in1(N__46729),
            .in2(N__42006),
            .in3(N__46831),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_6_f0_0_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_17_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_17_19_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_17_19_7  (
            .in0(N__46834),
            .in1(N__41645),
            .in2(N__41598),
            .in3(N__41494),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45966),
            .ce(N__46577),
            .sr(N__45500));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_17_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_17_20_0 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_17_20_0  (
            .in0(N__46844),
            .in1(N__46717),
            .in2(N__41594),
            .in3(N__41493),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45960),
            .ce(N__46581),
            .sr(N__45509));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_17_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_17_20_1 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_17_20_1  (
            .in0(N__41492),
            .in1(N__41374),
            .in2(N__46734),
            .in3(N__46846),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45960),
            .ce(N__46581),
            .sr(N__45509));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6_19_LC_17_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6_19_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6_19_LC_17_20_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6_19_LC_17_20_4  (
            .in0(N__41252),
            .in1(N__42089),
            .in2(N__41328),
            .in3(N__42101),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_6_f0_i_a2_0_6Z0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_17_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_17_20_7 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_17_20_7  (
            .in0(N__46716),
            .in1(N__41866),
            .in2(_gnd_net_),
            .in3(N__46845),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45960),
            .ce(N__46581),
            .sr(N__45509));
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_17_21_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_17_21_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_6_LC_17_21_1 .LUT_INIT=16'b1110101011111011;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_6_LC_17_21_1  (
            .in0(N__46460),
            .in1(N__46253),
            .in2(N__41292),
            .in3(N__42294),
            .lcout(measured_delay_hc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45955),
            .ce(),
            .sr(N__45516));
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_17_21_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_17_21_2 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_29_LC_17_21_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_29_LC_17_21_2  (
            .in0(N__46251),
            .in1(_gnd_net_),
            .in2(N__46493),
            .in3(N__41253),
            .lcout(measured_delay_hc_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45955),
            .ce(),
            .sr(N__45516));
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_17_21_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_17_21_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_27_LC_17_21_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_27_LC_17_21_3  (
            .in0(N__42102),
            .in1(N__46452),
            .in2(_gnd_net_),
            .in3(N__46249),
            .lcout(measured_delay_hc_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45955),
            .ce(),
            .sr(N__45516));
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_17_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_17_21_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_28_LC_17_21_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_28_LC_17_21_4  (
            .in0(N__46250),
            .in1(_gnd_net_),
            .in2(N__46492),
            .in3(N__42090),
            .lcout(measured_delay_hc_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45955),
            .ce(),
            .sr(N__45516));
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_17_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_17_21_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_31_LC_17_21_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_31_LC_17_21_5  (
            .in0(N__46713),
            .in1(N__46459),
            .in2(_gnd_net_),
            .in3(N__46252),
            .lcout(measured_delay_hc_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45955),
            .ce(),
            .sr(N__45516));
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_17_21_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_17_21_7 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_0_LC_17_21_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_0_LC_17_21_7  (
            .in0(N__42066),
            .in1(N__46451),
            .in2(_gnd_net_),
            .in3(N__46248),
            .lcout(measured_delay_hc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45955),
            .ce(),
            .sr(N__45516));
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_17_22_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_17_22_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_19_LC_17_22_1 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_19_LC_17_22_1  (
            .in0(N__46176),
            .in1(N__42045),
            .in2(N__46449),
            .in3(N__41997),
            .lcout(measured_delay_hc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45952),
            .ce(),
            .sr(N__45525));
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_17_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_17_22_4 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_16_LC_17_22_4 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_16_LC_17_22_4  (
            .in0(N__41961),
            .in1(N__46387),
            .in2(N__46994),
            .in3(N__46174),
            .lcout(measured_delay_hc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45952),
            .ce(),
            .sr(N__45525));
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_17_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_17_22_5 .SEQ_MODE=4'b1001;
    defparam \delay_measurement_inst.delay_hc_reg_1_LC_17_22_5 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_1_LC_17_22_5  (
            .in0(N__46177),
            .in1(N__42423),
            .in2(N__46450),
            .in3(N__41921),
            .lcout(measured_delay_hc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45952),
            .ce(),
            .sr(N__45525));
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_17_22_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_17_22_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_18_LC_17_22_6 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_18_LC_17_22_6  (
            .in0(N__41858),
            .in1(N__46388),
            .in2(N__41895),
            .in3(N__46175),
            .lcout(measured_delay_hc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45952),
            .ce(),
            .sr(N__45525));
    defparam reset_ibuf_gb_io_RNI79U7_LC_17_23_0.C_ON=1'b0;
    defparam reset_ibuf_gb_io_RNI79U7_LC_17_23_0.SEQ_MODE=4'b0000;
    defparam reset_ibuf_gb_io_RNI79U7_LC_17_23_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 reset_ibuf_gb_io_RNI79U7_LC_17_23_0 (
            .in0(N__45619),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(red_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_17_23_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_17_23_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJG9N1_1_LC_17_23_1  (
            .in0(N__42422),
            .in1(N__46304),
            .in2(N__42405),
            .in3(N__42371),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_reg3_i_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_17_24_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_17_24_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_17_24_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_RNO_0_6_LC_17_24_7  (
            .in0(N__42339),
            .in1(N__42317),
            .in2(_gnd_net_),
            .in3(N__42305),
            .lcout(\delay_measurement_inst.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_17_25_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_17_25_1 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_15_LC_17_25_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_15_LC_17_25_1  (
            .in0(N__42285),
            .in1(N__46352),
            .in2(N__42256),
            .in3(N__46254),
            .lcout(measured_delay_hc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45944),
            .ce(),
            .sr(N__45547));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_9_0 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_9_0  (
            .in0(N__42617),
            .in1(N__42938),
            .in2(N__42213),
            .in3(N__42814),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46054),
            .ce(),
            .sr(N__45442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_9_1 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_9_1  (
            .in0(N__42813),
            .in1(N__42619),
            .in2(N__42959),
            .in3(N__42168),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46054),
            .ce(),
            .sr(N__45442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_9_2 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_9_2  (
            .in0(N__42618),
            .in1(N__42939),
            .in2(N__42132),
            .in3(N__42815),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46054),
            .ce(),
            .sr(N__45442));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_18_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_18_9_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_LC_18_9_4  (
            .in0(N__43953),
            .in1(N__44221),
            .in2(_gnd_net_),
            .in3(N__47069),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_9_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_9_5  (
            .in0(N__44473),
            .in1(N__44666),
            .in2(N__42105),
            .in3(N__44357),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46054),
            .ce(),
            .sr(N__45442));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_9_7 .LUT_INIT=16'b1111100100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_9_7  (
            .in0(N__44472),
            .in1(N__44667),
            .in2(N__44358),
            .in3(N__44010),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46054),
            .ce(),
            .sr(N__45442));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__43880),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46046),
            .ce(N__43828),
            .sr(N__45445));
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_18_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_18_11_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_17_LC_18_11_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_17_LC_18_11_5  (
            .in0(N__43672),
            .in1(N__43805),
            .in2(_gnd_net_),
            .in3(N__43730),
            .lcout(measured_delay_tr_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46038),
            .ce(N__43515),
            .sr(N__45448));
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_18_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_tr_reg_esr_18_LC_18_11_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_reg_esr_18_LC_18_11_6  (
            .in0(N__43731),
            .in1(N__43673),
            .in2(_gnd_net_),
            .in3(N__43581),
            .lcout(measured_delay_tr_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46038),
            .ce(N__43515),
            .sr(N__45448));
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.stoper_state_1_LC_18_12_1 .LUT_INIT=16'b0100000001001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.stoper_state_1_LC_18_12_1  (
            .in0(N__43450),
            .in1(N__43330),
            .in2(N__43031),
            .in3(N__43176),
            .lcout(\phase_controller_inst1.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__42510),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.stoper_state_1_LC_18_12_3 .LUT_INIT=16'b0000100001011000;
    LogicCell40 \phase_controller_inst1.stoper_tr.stoper_state_1_LC_18_12_3  (
            .in0(N__42540),
            .in1(N__42943),
            .in2(N__42819),
            .in3(N__42680),
            .lcout(\phase_controller_inst1.stoper_tr.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__42510),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_18_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_0_LC_18_12_4 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_0_LC_18_12_4  (
            .in0(N__44444),
            .in1(N__44653),
            .in2(N__44340),
            .in3(N__47061),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__42510),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_18_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_18_12_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_1_LC_18_12_5 .LUT_INIT=16'b0001000111000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_1_LC_18_12_5  (
            .in0(N__47062),
            .in1(N__44445),
            .in2(N__44665),
            .in3(N__44298),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__46027),
            .ce(N__42510),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__43945),
            .in2(_gnd_net_),
            .in3(N__47059),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_18_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_18_12_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2P_LC_18_12_7  (
            .in0(N__47060),
            .in1(_gnd_net_),
            .in2(N__43952),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_RNIUO2PZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0_0_c_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__43923),
            .in2(N__44229),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_18_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_2_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__44184),
            .in2(_gnd_net_),
            .in3(N__43917),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_18_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_18_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_3_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__43914),
            .in2(N__44163),
            .in3(N__43908),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_18_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_18_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_4_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__44115),
            .in2(_gnd_net_),
            .in3(N__43905),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_18_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_18_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_5_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__44904),
            .in2(_gnd_net_),
            .in3(N__43902),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_18_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_18_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_6_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__44883),
            .in2(_gnd_net_),
            .in3(N__43899),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_18_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_18_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_7_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__44853),
            .in2(_gnd_net_),
            .in3(N__43887),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_18_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_18_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_8_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__44814),
            .in2(_gnd_net_),
            .in3(N__43884),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_18_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_18_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_9_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__44774),
            .in2(_gnd_net_),
            .in3(N__44013),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_9 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_18_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_18_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_10_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__44744),
            .in2(_gnd_net_),
            .in3(N__44001),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_18_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_18_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_11_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__44708),
            .in2(_gnd_net_),
            .in3(N__43992),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_18_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_18_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_12_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__45150),
            .in2(_gnd_net_),
            .in3(N__43989),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_18_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_18_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_13_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__45126),
            .in2(_gnd_net_),
            .in3(N__43977),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_18_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_18_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_14_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__45077),
            .in2(_gnd_net_),
            .in3(N__43974),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_18_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_18_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_15_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__45032),
            .in2(_gnd_net_),
            .in3(N__43965),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_18_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_18_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_16_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__45008),
            .in2(_gnd_net_),
            .in3(N__43956),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_18_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_18_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_17_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__44987),
            .in2(_gnd_net_),
            .in3(N__44088),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_17 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_18_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_18_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_18_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__44957),
            .in2(_gnd_net_),
            .in3(N__44079),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_18_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_18_15_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_19_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__44936),
            .in2(_gnd_net_),
            .in3(N__44076),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_RNO_0_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_18_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_18_15_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.stoper_state_RNI0RST_0_LC_18_15_4  (
            .in0(N__44560),
            .in1(N__44433),
            .in2(_gnd_net_),
            .in3(N__44302),
            .lcout(\phase_controller_inst2.stoper_hc.stoper_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_16_0 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_16_0  (
            .in0(N__44346),
            .in1(N__44646),
            .in2(N__44508),
            .in3(N__44067),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_16_1 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_16_1  (
            .in0(N__44645),
            .in1(N__44492),
            .in2(N__44058),
            .in3(N__44352),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_16_2 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_16_2  (
            .in0(N__44348),
            .in1(N__44648),
            .in2(N__44510),
            .in3(N__44046),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_16_3 .LUT_INIT=16'b1010101010000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_16_3  (
            .in0(N__44037),
            .in1(N__44489),
            .in2(N__44664),
            .in3(N__44353),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_16_4 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_16_4  (
            .in0(N__44347),
            .in1(N__44647),
            .in2(N__44509),
            .in3(N__44028),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_16_5 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_16_5  (
            .in0(N__44643),
            .in1(N__44490),
            .in2(N__44688),
            .in3(N__44350),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_16_6 .LUT_INIT=16'b1110101100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_16_6  (
            .in0(N__44349),
            .in1(N__44649),
            .in2(N__44511),
            .in3(N__44676),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_16_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_16_7  (
            .in0(N__44644),
            .in1(N__44491),
            .in2(N__44373),
            .in3(N__44351),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45992),
            .ce(),
            .sr(N__45479));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_18_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_18_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_18_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_18_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1_c_inv_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__44202),
            .in2(N__44238),
            .in3(N__44228),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_18_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_18_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2_c_inv_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__44169),
            .in2(N__44196),
            .in3(N__44180),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_18_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_18_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3_c_inv_LC_18_17_3  (
            .in0(N__44156),
            .in1(N__44130),
            .in2(N__44145),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_18_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_18_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4_c_inv_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__44100),
            .in2(N__44124),
            .in3(N__44111),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_18_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_18_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5_c_inv_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__44889),
            .in2(N__44916),
            .in3(N__44900),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_18_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_18_17_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6_c_inv_LC_18_17_6  (
            .in0(N__44879),
            .in1(N__44859),
            .in2(N__44868),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_18_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_18_17_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7_c_inv_LC_18_17_7  (
            .in0(N__44849),
            .in1(N__44826),
            .in2(N__44838),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_18_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_18_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8_c_inv_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__44820),
            .in2(N__44796),
            .in3(N__44813),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_18_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_18_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9_c_inv_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__44760),
            .in2(N__44787),
            .in3(N__44775),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_18_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_18_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10_c_inv_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__44727),
            .in2(N__44754),
            .in3(N__44745),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_18_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_18_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11_c_inv_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__44694),
            .in2(N__44721),
            .in3(N__44712),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_18_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_18_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12_c_inv_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__45132),
            .in2(N__45159),
            .in3(N__45149),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_18_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_18_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13_c_inv_LC_18_18_5  (
            .in0(N__45122),
            .in1(N__45096),
            .in2(N__45108),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_18_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_18_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14_c_inv_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__45090),
            .in2(N__45057),
            .in3(N__45078),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_18_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_18_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15_c_inv_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__45018),
            .in2(N__45048),
            .in3(N__45036),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_18_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_18_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16_c_inv_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__44994),
            .in2(N__46956),
            .in3(N__45012),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_16 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_18_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_18_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17_c_inv_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__44973),
            .in2(N__46593),
            .in3(N__44988),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_18_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_18_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18_c_inv_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__44943),
            .in2(N__44967),
            .in3(N__44958),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_18_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_18_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_c_inv_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__44922),
            .in2(N__47004),
            .in3(N__44937),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_LUT4_0_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47073),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_18_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_18_20_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__46712),
            .in2(_gnd_net_),
            .in3(N__47028),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45967),
            .ce(N__46580),
            .sr(N__45501));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_21_6 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_18_21_6  (
            .in0(N__46714),
            .in1(N__46984),
            .in2(_gnd_net_),
            .in3(N__46917),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45961),
            .ce(N__46578),
            .sr(N__45510));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_21_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_18_21_7  (
            .in0(N__46916),
            .in1(N__46715),
            .in2(_gnd_net_),
            .in3(N__46647),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45961),
            .ce(N__46578),
            .sr(N__45510));
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_18_22_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_25_LC_18_22_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_25_LC_18_22_3  (
            .in0(N__46514),
            .in1(N__46482),
            .in2(_gnd_net_),
            .in3(N__46276),
            .lcout(measured_delay_hc_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45956),
            .ce(),
            .sr(N__45517));
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_18_22_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_18_22_5 .SEQ_MODE=4'b1000;
    defparam \delay_measurement_inst.delay_hc_reg_2_LC_18_22_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_reg_2_LC_18_22_5  (
            .in0(N__46112),
            .in1(N__46483),
            .in2(N__46311),
            .in3(N__46277),
            .lcout(measured_delay_hc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__45956),
            .ce(),
            .sr(N__45517));
endmodule // MAIN
